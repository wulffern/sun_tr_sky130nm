magic
tech sky130B
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 1260 1056
<< locali >>
rect 168 58 396 118
rect 168 938 396 998
rect 168 58 228 998
rect 396 410 564 470
rect 396 586 564 646
rect 564 410 624 646
rect 798 146 858 734
rect 366 410 426 646
rect 1152 132 1368 220
rect 288 410 504 470
rect 720 146 936 206
rect 288 58 504 118
use SUNTR_PCHDLCM M0
transform 1 0 0 0 1 0
box 0 0 1260 528
use SUNTR_PCHDLCM M1
transform 1 0 0 0 1 528
box 0 528 1260 1056
<< labels >>
flabel locali s 1152 132 1368 220 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel locali s 288 410 504 470 0 FreeSans 400 0 0 0 D
port 1 nsew
flabel locali s 720 146 936 206 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 288 58 504 118 0 FreeSans 400 0 0 0 S
port 3 nsew
<< end >>
