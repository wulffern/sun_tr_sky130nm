magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 2672 4236
<< locali >>
rect 16 16 2656 128
rect 128 16 2544 128
rect 16 16 2656 128
rect 128 4108 2544 4220
rect 16 4108 2656 4220
rect 16 128 128 4108
rect 16 16 128 4220
rect 2544 128 2656 4108
rect 2544 16 2656 4220
rect 16 16 2656 128
rect 1480 3438 2056 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 176 32 256 112
rect 256 32 336 112
rect 336 32 416 112
rect 416 32 496 112
rect 496 32 576 112
rect 576 32 656 112
rect 656 32 736 112
rect 736 32 816 112
rect 816 32 896 112
rect 896 32 976 112
rect 976 32 1056 112
rect 1056 32 1136 112
rect 1136 32 1216 112
rect 1216 32 1296 112
rect 1296 32 1376 112
rect 1376 32 1456 112
rect 1456 32 1536 112
rect 1536 32 1616 112
rect 1616 32 1696 112
rect 1696 32 1776 112
rect 1776 32 1856 112
rect 1856 32 1936 112
rect 1936 32 2016 112
rect 2016 32 2096 112
rect 2096 32 2176 112
rect 2176 32 2256 112
rect 2256 32 2336 112
rect 2336 32 2416 112
rect 2416 32 2496 112
rect 176 4124 256 4204
rect 256 4124 336 4204
rect 336 4124 416 4204
rect 416 4124 496 4204
rect 496 4124 576 4204
rect 576 4124 656 4204
rect 656 4124 736 4204
rect 736 4124 816 4204
rect 816 4124 896 4204
rect 896 4124 976 4204
rect 976 4124 1056 4204
rect 1056 4124 1136 4204
rect 1136 4124 1216 4204
rect 1216 4124 1296 4204
rect 1296 4124 1376 4204
rect 1376 4124 1456 4204
rect 1456 4124 1536 4204
rect 1536 4124 1616 4204
rect 1616 4124 1696 4204
rect 1696 4124 1776 4204
rect 1776 4124 1856 4204
rect 1856 4124 1936 4204
rect 1936 4124 2016 4204
rect 2016 4124 2096 4204
rect 2096 4124 2176 4204
rect 2176 4124 2256 4204
rect 2256 4124 2336 4204
rect 2336 4124 2416 4204
rect 2416 4124 2496 4204
rect 32 158 112 238
rect 32 238 112 318
rect 32 318 112 398
rect 32 398 112 478
rect 32 478 112 558
rect 32 558 112 638
rect 32 638 112 718
rect 32 718 112 798
rect 32 798 112 878
rect 32 878 112 958
rect 32 958 112 1038
rect 32 1038 112 1118
rect 32 1118 112 1198
rect 32 1198 112 1278
rect 32 1278 112 1358
rect 32 1358 112 1438
rect 32 1438 112 1518
rect 32 1518 112 1598
rect 32 1598 112 1678
rect 32 1678 112 1758
rect 32 1758 112 1838
rect 32 1838 112 1918
rect 32 1918 112 1998
rect 32 1998 112 2078
rect 32 2078 112 2158
rect 32 2158 112 2238
rect 32 2238 112 2318
rect 32 2318 112 2398
rect 32 2398 112 2478
rect 32 2478 112 2558
rect 32 2558 112 2638
rect 32 2638 112 2718
rect 32 2718 112 2798
rect 32 2798 112 2878
rect 32 2878 112 2958
rect 32 2958 112 3038
rect 32 3038 112 3118
rect 32 3118 112 3198
rect 32 3198 112 3278
rect 32 3278 112 3358
rect 32 3358 112 3438
rect 32 3438 112 3518
rect 32 3518 112 3598
rect 32 3598 112 3678
rect 32 3678 112 3758
rect 32 3758 112 3838
rect 32 3838 112 3918
rect 32 3918 112 3998
rect 32 3998 112 4078
rect 2560 158 2640 238
rect 2560 238 2640 318
rect 2560 318 2640 398
rect 2560 398 2640 478
rect 2560 478 2640 558
rect 2560 558 2640 638
rect 2560 638 2640 718
rect 2560 718 2640 798
rect 2560 798 2640 878
rect 2560 878 2640 958
rect 2560 958 2640 1038
rect 2560 1038 2640 1118
rect 2560 1118 2640 1198
rect 2560 1198 2640 1278
rect 2560 1278 2640 1358
rect 2560 1358 2640 1438
rect 2560 1438 2640 1518
rect 2560 1518 2640 1598
rect 2560 1598 2640 1678
rect 2560 1678 2640 1758
rect 2560 1758 2640 1838
rect 2560 1838 2640 1918
rect 2560 1918 2640 1998
rect 2560 1998 2640 2078
rect 2560 2078 2640 2158
rect 2560 2158 2640 2238
rect 2560 2238 2640 2318
rect 2560 2318 2640 2398
rect 2560 2398 2640 2478
rect 2560 2478 2640 2558
rect 2560 2558 2640 2638
rect 2560 2638 2640 2718
rect 2560 2718 2640 2798
rect 2560 2798 2640 2878
rect 2560 2878 2640 2958
rect 2560 2958 2640 3038
rect 2560 3038 2640 3118
rect 2560 3118 2640 3198
rect 2560 3198 2640 3278
rect 2560 3278 2640 3358
rect 2560 3358 2640 3438
rect 2560 3438 2640 3518
rect 2560 3518 2640 3598
rect 2560 3598 2640 3678
rect 2560 3678 2640 3758
rect 2560 3758 2640 3838
rect 2560 3838 2640 3918
rect 2560 3918 2640 3998
rect 2560 3998 2640 4078
<< ptap >>
rect 0 0 2672 144
rect 0 4092 2672 4236
rect 0 0 144 4236
rect 2528 0 2672 4236
use SUNTR_RES2 XA1 
transform 1 0 688 0 1 688
box 688 688 1984 3548
<< labels >>
flabel locali s 16 16 2656 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 1480 3438 2056 3658 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2672 4236
<< end >>
