magic
tech sky130B
timestamp 1728046668
<< psubdiff >>
rect 0 2102 2632 2118
rect 0 2062 76 2102
rect 2556 2062 2632 2102
rect 0 2046 2632 2062
rect 0 2039 72 2046
rect 0 79 16 2039
rect 56 79 72 2039
rect 0 72 72 79
rect 2560 2039 2632 2046
rect 2560 79 2576 2039
rect 2616 79 2632 2039
rect 2560 72 2632 79
rect 0 56 2632 72
rect 0 16 76 56
rect 2556 16 2632 56
rect 0 0 2632 16
<< psubdiffcont >>
rect 76 2062 2556 2102
rect 16 79 56 2039
rect 2576 79 2616 2039
rect 76 16 2556 56
<< locali >>
rect 8 2102 2624 2110
rect 8 2062 76 2102
rect 2556 2062 2624 2102
rect 8 2054 2624 2062
rect 8 2039 64 2054
rect 8 79 16 2039
rect 56 79 64 2039
rect 2568 2039 2624 2054
rect 308 1719 596 1829
rect 2036 1719 2324 1829
rect 8 64 64 79
rect 2568 79 2576 2039
rect 2616 79 2624 2039
rect 2568 64 2624 79
rect 8 56 2624 64
rect 8 16 76 56
rect 2556 16 2624 56
rect 8 8 2624 16
use SUNTR_RES8  XA1
timestamp 1709161200
transform 1 0 344 0 1 344
box -36 -55 1980 1485
<< labels >>
flabel locali s 8 8 2624 64 0 FreeSans 200 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 2036 1719 2324 1829 0 FreeSans 200 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 308 1719 596 1829 0 FreeSans 200 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2632 2118
<< end >>
