* NGSPICE file created from SUNTR_NCHL.ext - technology: sky130B

.subckt SUNTR_NCHL D G S B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=5.184e+11p pd=3.12e+06u as=5.184e+11p ps=3.12e+06u w=1.08e+06u l=360000u
C0 a_324_n36# B 0.43fF $ **FLOATING
C1 a_324_492# B 0.43fF $ **FLOATING
.ends
