*idgm_lvt

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../design/SUN_TR_SKY130NM.spice

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
*.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

.param dv = 1n

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD 0 dc 1.8
INN N1_REF 0 dc {dv}
VREF N1_REF VDD dc 0.5

BINN 0 N1 i=i(VREF) tc1=0

E0 EN0 VDD N1 VDD 1
E1 EN1 VDD N1 VDD 1
E2 EN2 VDD N1 VDD 1
VD1 N2 N1 dc {dv}
VD2 EN3 EN2 dc {dv}

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
XM1 N1 N1 VDD VDD SUNTR_PCHDL
XM2 EN0 N1 VDD VDD SUNTR_PCHDL
XM3 EN1 N2 VDD VDD SUNTR_PCHDL
XM4 EN3 N1 VDD VDD SUNTR_PCHDL

B1 gm 0 v=(i(E0) - i(E1))/{dv}
B2 idsq 0 v=i(INN)/3
B3 gmid 0 v=v(gm)/i(inn)
B4 vgs 0 v=v(vdd)-v(n1)
B5 rds 0 v={dv}/(i(E0) - i(E2))
B6 gmrds 0 v=v(gm)*v(rds)
B7 gmrds_db 0 v=20*log10(abs(v(gm)*v(rds)))

*.save @XM1.XMM1M1[gm]

.probe i(inn) i(e0) i(e1) v(n1) v(gm) v(EN1) v(EN0) v(idsq) v(gmid) v(vgs)
*----------------------------------------------------------------
* Control
*----------------------------------------------------------------
.control
unset askquit
dc inn 1n 100u 100n
write
quit
.endc
.end
