* NGSPICE file created from SUNTR_CAP_20.ext - technology: sky130B

.subckt SUNTR_CAP_20 A B
R0 A m3_5076_132# sky130_fd_pr__res_generic_m3 w=440000u l=360000u
R1 m3_252_308# B sky130_fd_pr__res_generic_m3 w=440000u l=360000u
C0 A B 36.69fF
C1 B 0 8.91fF
C2 A 0 8.87fF
.ends
