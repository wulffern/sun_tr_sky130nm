magic
tech sky130B
magscale 1 2
timestamp 1709161200
<< checkpaint >>
rect 0 0 8720 4236
<< locali >>
rect 16 16 8704 128
rect 128 16 8592 128
rect 16 16 8704 128
rect 128 4108 8592 4220
rect 16 4108 8704 4220
rect 16 128 128 4108
rect 16 16 128 4220
rect 8592 128 8704 4108
rect 8592 16 8704 4220
rect 16 16 8704 128
rect 7528 3438 8104 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 160 32 240 112
rect 240 32 320 112
rect 320 32 400 112
rect 400 32 480 112
rect 480 32 560 112
rect 560 32 640 112
rect 640 32 720 112
rect 720 32 800 112
rect 800 32 880 112
rect 880 32 960 112
rect 960 32 1040 112
rect 1040 32 1120 112
rect 1120 32 1200 112
rect 1200 32 1280 112
rect 1280 32 1360 112
rect 1360 32 1440 112
rect 1440 32 1520 112
rect 1520 32 1600 112
rect 1600 32 1680 112
rect 1680 32 1760 112
rect 1760 32 1840 112
rect 1840 32 1920 112
rect 1920 32 2000 112
rect 2000 32 2080 112
rect 2080 32 2160 112
rect 2160 32 2240 112
rect 2240 32 2320 112
rect 2320 32 2400 112
rect 2400 32 2480 112
rect 2480 32 2560 112
rect 2560 32 2640 112
rect 2640 32 2720 112
rect 2720 32 2800 112
rect 2800 32 2880 112
rect 2880 32 2960 112
rect 2960 32 3040 112
rect 3040 32 3120 112
rect 3120 32 3200 112
rect 3200 32 3280 112
rect 3280 32 3360 112
rect 3360 32 3440 112
rect 3440 32 3520 112
rect 3520 32 3600 112
rect 3600 32 3680 112
rect 3680 32 3760 112
rect 3760 32 3840 112
rect 3840 32 3920 112
rect 3920 32 4000 112
rect 4000 32 4080 112
rect 4080 32 4160 112
rect 4160 32 4240 112
rect 4240 32 4320 112
rect 4320 32 4400 112
rect 4400 32 4480 112
rect 4480 32 4560 112
rect 4560 32 4640 112
rect 4640 32 4720 112
rect 4720 32 4800 112
rect 4800 32 4880 112
rect 4880 32 4960 112
rect 4960 32 5040 112
rect 5040 32 5120 112
rect 5120 32 5200 112
rect 5200 32 5280 112
rect 5280 32 5360 112
rect 5360 32 5440 112
rect 5440 32 5520 112
rect 5520 32 5600 112
rect 5600 32 5680 112
rect 5680 32 5760 112
rect 5760 32 5840 112
rect 5840 32 5920 112
rect 5920 32 6000 112
rect 6000 32 6080 112
rect 6080 32 6160 112
rect 6160 32 6240 112
rect 6240 32 6320 112
rect 6320 32 6400 112
rect 6400 32 6480 112
rect 6480 32 6560 112
rect 6560 32 6640 112
rect 6640 32 6720 112
rect 6720 32 6800 112
rect 6800 32 6880 112
rect 6880 32 6960 112
rect 6960 32 7040 112
rect 7040 32 7120 112
rect 7120 32 7200 112
rect 7200 32 7280 112
rect 7280 32 7360 112
rect 7360 32 7440 112
rect 7440 32 7520 112
rect 7520 32 7600 112
rect 7600 32 7680 112
rect 7680 32 7760 112
rect 7760 32 7840 112
rect 7840 32 7920 112
rect 7920 32 8000 112
rect 8000 32 8080 112
rect 8080 32 8160 112
rect 8160 32 8240 112
rect 8240 32 8320 112
rect 8320 32 8400 112
rect 8400 32 8480 112
rect 8480 32 8560 112
rect 160 4124 240 4204
rect 240 4124 320 4204
rect 320 4124 400 4204
rect 400 4124 480 4204
rect 480 4124 560 4204
rect 560 4124 640 4204
rect 640 4124 720 4204
rect 720 4124 800 4204
rect 800 4124 880 4204
rect 880 4124 960 4204
rect 960 4124 1040 4204
rect 1040 4124 1120 4204
rect 1120 4124 1200 4204
rect 1200 4124 1280 4204
rect 1280 4124 1360 4204
rect 1360 4124 1440 4204
rect 1440 4124 1520 4204
rect 1520 4124 1600 4204
rect 1600 4124 1680 4204
rect 1680 4124 1760 4204
rect 1760 4124 1840 4204
rect 1840 4124 1920 4204
rect 1920 4124 2000 4204
rect 2000 4124 2080 4204
rect 2080 4124 2160 4204
rect 2160 4124 2240 4204
rect 2240 4124 2320 4204
rect 2320 4124 2400 4204
rect 2400 4124 2480 4204
rect 2480 4124 2560 4204
rect 2560 4124 2640 4204
rect 2640 4124 2720 4204
rect 2720 4124 2800 4204
rect 2800 4124 2880 4204
rect 2880 4124 2960 4204
rect 2960 4124 3040 4204
rect 3040 4124 3120 4204
rect 3120 4124 3200 4204
rect 3200 4124 3280 4204
rect 3280 4124 3360 4204
rect 3360 4124 3440 4204
rect 3440 4124 3520 4204
rect 3520 4124 3600 4204
rect 3600 4124 3680 4204
rect 3680 4124 3760 4204
rect 3760 4124 3840 4204
rect 3840 4124 3920 4204
rect 3920 4124 4000 4204
rect 4000 4124 4080 4204
rect 4080 4124 4160 4204
rect 4160 4124 4240 4204
rect 4240 4124 4320 4204
rect 4320 4124 4400 4204
rect 4400 4124 4480 4204
rect 4480 4124 4560 4204
rect 4560 4124 4640 4204
rect 4640 4124 4720 4204
rect 4720 4124 4800 4204
rect 4800 4124 4880 4204
rect 4880 4124 4960 4204
rect 4960 4124 5040 4204
rect 5040 4124 5120 4204
rect 5120 4124 5200 4204
rect 5200 4124 5280 4204
rect 5280 4124 5360 4204
rect 5360 4124 5440 4204
rect 5440 4124 5520 4204
rect 5520 4124 5600 4204
rect 5600 4124 5680 4204
rect 5680 4124 5760 4204
rect 5760 4124 5840 4204
rect 5840 4124 5920 4204
rect 5920 4124 6000 4204
rect 6000 4124 6080 4204
rect 6080 4124 6160 4204
rect 6160 4124 6240 4204
rect 6240 4124 6320 4204
rect 6320 4124 6400 4204
rect 6400 4124 6480 4204
rect 6480 4124 6560 4204
rect 6560 4124 6640 4204
rect 6640 4124 6720 4204
rect 6720 4124 6800 4204
rect 6800 4124 6880 4204
rect 6880 4124 6960 4204
rect 6960 4124 7040 4204
rect 7040 4124 7120 4204
rect 7120 4124 7200 4204
rect 7200 4124 7280 4204
rect 7280 4124 7360 4204
rect 7360 4124 7440 4204
rect 7440 4124 7520 4204
rect 7520 4124 7600 4204
rect 7600 4124 7680 4204
rect 7680 4124 7760 4204
rect 7760 4124 7840 4204
rect 7840 4124 7920 4204
rect 7920 4124 8000 4204
rect 8000 4124 8080 4204
rect 8080 4124 8160 4204
rect 8160 4124 8240 4204
rect 8240 4124 8320 4204
rect 8320 4124 8400 4204
rect 8400 4124 8480 4204
rect 8480 4124 8560 4204
rect 32 158 112 238
rect 32 238 112 318
rect 32 318 112 398
rect 32 398 112 478
rect 32 478 112 558
rect 32 558 112 638
rect 32 638 112 718
rect 32 718 112 798
rect 32 798 112 878
rect 32 878 112 958
rect 32 958 112 1038
rect 32 1038 112 1118
rect 32 1118 112 1198
rect 32 1198 112 1278
rect 32 1278 112 1358
rect 32 1358 112 1438
rect 32 1438 112 1518
rect 32 1518 112 1598
rect 32 1598 112 1678
rect 32 1678 112 1758
rect 32 1758 112 1838
rect 32 1838 112 1918
rect 32 1918 112 1998
rect 32 1998 112 2078
rect 32 2078 112 2158
rect 32 2158 112 2238
rect 32 2238 112 2318
rect 32 2318 112 2398
rect 32 2398 112 2478
rect 32 2478 112 2558
rect 32 2558 112 2638
rect 32 2638 112 2718
rect 32 2718 112 2798
rect 32 2798 112 2878
rect 32 2878 112 2958
rect 32 2958 112 3038
rect 32 3038 112 3118
rect 32 3118 112 3198
rect 32 3198 112 3278
rect 32 3278 112 3358
rect 32 3358 112 3438
rect 32 3438 112 3518
rect 32 3518 112 3598
rect 32 3598 112 3678
rect 32 3678 112 3758
rect 32 3758 112 3838
rect 32 3838 112 3918
rect 32 3918 112 3998
rect 32 3998 112 4078
rect 8608 158 8688 238
rect 8608 238 8688 318
rect 8608 318 8688 398
rect 8608 398 8688 478
rect 8608 478 8688 558
rect 8608 558 8688 638
rect 8608 638 8688 718
rect 8608 718 8688 798
rect 8608 798 8688 878
rect 8608 878 8688 958
rect 8608 958 8688 1038
rect 8608 1038 8688 1118
rect 8608 1118 8688 1198
rect 8608 1198 8688 1278
rect 8608 1278 8688 1358
rect 8608 1358 8688 1438
rect 8608 1438 8688 1518
rect 8608 1518 8688 1598
rect 8608 1598 8688 1678
rect 8608 1678 8688 1758
rect 8608 1758 8688 1838
rect 8608 1838 8688 1918
rect 8608 1918 8688 1998
rect 8608 1998 8688 2078
rect 8608 2078 8688 2158
rect 8608 2158 8688 2238
rect 8608 2238 8688 2318
rect 8608 2318 8688 2398
rect 8608 2398 8688 2478
rect 8608 2478 8688 2558
rect 8608 2558 8688 2638
rect 8608 2638 8688 2718
rect 8608 2718 8688 2798
rect 8608 2798 8688 2878
rect 8608 2878 8688 2958
rect 8608 2958 8688 3038
rect 8608 3038 8688 3118
rect 8608 3118 8688 3198
rect 8608 3198 8688 3278
rect 8608 3278 8688 3358
rect 8608 3358 8688 3438
rect 8608 3438 8688 3518
rect 8608 3518 8688 3598
rect 8608 3598 8688 3678
rect 8608 3678 8688 3758
rect 8608 3758 8688 3838
rect 8608 3838 8688 3918
rect 8608 3918 8688 3998
rect 8608 3998 8688 4078
<< ptap >>
rect 0 0 8720 144
rect 0 4092 8720 4236
rect 0 0 144 4236
rect 8576 0 8720 4236
use SUNTR_RES16 XA1 
transform 1 0 688 0 1 688
box 688 688 8032 3548
<< labels >>
flabel locali s 16 16 8704 128 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 7528 3438 8104 3658 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 8720 4236
<< end >>
