*idgm_lvt

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../design/SUN_TR_SKY130NM.spice

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VSS VSS 0 dc 0
INN 0 N1_REF dc 1u
VREF N1_REF 0 dc 0.5

BINN 0 N1 i=i(VREF) tc1=0

E0 EN0 0 N1 0 1
E1 EN1 0 N1 0 1
E2 EN2 0 N1 0 1
VD1 N2 N1 dc 1u
VD2 EN3 EN2 dc 1m

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
XM1 N1 N1 VSS VSS SUNTR_NCHDL
XM2 EN0 N1 VSS VSS SUNTR_NCHDL
XM3 EN1 N2 VSS VSS SUNTR_NCHDL
XM4 EN3 N1 VSS VSS SUNTR_NCHDL

B1 gm 0 v=(i(E0) - i(E1))/1u
B2 idsq 0 v=i(INN)/3
B3 gmid 0 v=v(gm)/i(inn)
B4 rds 0 v=1m/(i(E0) - i(E2))
B5 gmrds 0 v=v(gm)*v(rds)
B6 gmrds_db 0 v=20*log10(abs(v(gm)*v(rds)))


.probe i(inn) i(e0) i(e1) v(n1) v(gm) v(EN1) v(EN0) v(idsq) v(gmid)
*----------------------------------------------------------------
* Control
*----------------------------------------------------------------
.control
unset askquit
dc inn 0.001u 100u 0.01u
write
quit
.endc
.end
