magic
tech sky130B
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 5264 4236
<< locali >>
rect 16 16 5248 128
rect 128 16 5136 128
rect 128 4108 5136 4220
rect 16 128 128 4108
rect 5136 128 5248 4108
rect 16 16 5248 128
rect 4072 3438 4648 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 152 32 232 112
rect 232 32 312 112
rect 312 32 392 112
rect 392 32 472 112
rect 472 32 552 112
rect 552 32 632 112
rect 632 32 712 112
rect 712 32 792 112
rect 792 32 872 112
rect 872 32 952 112
rect 952 32 1032 112
rect 1032 32 1112 112
rect 1112 32 1192 112
rect 1192 32 1272 112
rect 1272 32 1352 112
rect 1352 32 1432 112
rect 1432 32 1512 112
rect 1512 32 1592 112
rect 1592 32 1672 112
rect 1672 32 1752 112
rect 1752 32 1832 112
rect 1832 32 1912 112
rect 1912 32 1992 112
rect 1992 32 2072 112
rect 2072 32 2152 112
rect 2152 32 2232 112
rect 2232 32 2312 112
rect 2312 32 2392 112
rect 2392 32 2472 112
rect 2472 32 2552 112
rect 2552 32 2632 112
rect 2632 32 2712 112
rect 2712 32 2792 112
rect 2792 32 2872 112
rect 2872 32 2952 112
rect 2952 32 3032 112
rect 3032 32 3112 112
rect 3112 32 3192 112
rect 3192 32 3272 112
rect 3272 32 3352 112
rect 3352 32 3432 112
rect 3432 32 3512 112
rect 3512 32 3592 112
rect 3592 32 3672 112
rect 3672 32 3752 112
rect 3752 32 3832 112
rect 3832 32 3912 112
rect 3912 32 3992 112
rect 3992 32 4072 112
rect 4072 32 4152 112
rect 4152 32 4232 112
rect 4232 32 4312 112
rect 4312 32 4392 112
rect 4392 32 4472 112
rect 4472 32 4552 112
rect 4552 32 4632 112
rect 4632 32 4712 112
rect 4712 32 4792 112
rect 4792 32 4872 112
rect 4872 32 4952 112
rect 4952 32 5032 112
rect 5032 32 5112 112
rect 152 4124 232 4204
rect 232 4124 312 4204
rect 312 4124 392 4204
rect 392 4124 472 4204
rect 472 4124 552 4204
rect 552 4124 632 4204
rect 632 4124 712 4204
rect 712 4124 792 4204
rect 792 4124 872 4204
rect 872 4124 952 4204
rect 952 4124 1032 4204
rect 1032 4124 1112 4204
rect 1112 4124 1192 4204
rect 1192 4124 1272 4204
rect 1272 4124 1352 4204
rect 1352 4124 1432 4204
rect 1432 4124 1512 4204
rect 1512 4124 1592 4204
rect 1592 4124 1672 4204
rect 1672 4124 1752 4204
rect 1752 4124 1832 4204
rect 1832 4124 1912 4204
rect 1912 4124 1992 4204
rect 1992 4124 2072 4204
rect 2072 4124 2152 4204
rect 2152 4124 2232 4204
rect 2232 4124 2312 4204
rect 2312 4124 2392 4204
rect 2392 4124 2472 4204
rect 2472 4124 2552 4204
rect 2552 4124 2632 4204
rect 2632 4124 2712 4204
rect 2712 4124 2792 4204
rect 2792 4124 2872 4204
rect 2872 4124 2952 4204
rect 2952 4124 3032 4204
rect 3032 4124 3112 4204
rect 3112 4124 3192 4204
rect 3192 4124 3272 4204
rect 3272 4124 3352 4204
rect 3352 4124 3432 4204
rect 3432 4124 3512 4204
rect 3512 4124 3592 4204
rect 3592 4124 3672 4204
rect 3672 4124 3752 4204
rect 3752 4124 3832 4204
rect 3832 4124 3912 4204
rect 3912 4124 3992 4204
rect 3992 4124 4072 4204
rect 4072 4124 4152 4204
rect 4152 4124 4232 4204
rect 4232 4124 4312 4204
rect 4312 4124 4392 4204
rect 4392 4124 4472 4204
rect 4472 4124 4552 4204
rect 4552 4124 4632 4204
rect 4632 4124 4712 4204
rect 4712 4124 4792 4204
rect 4792 4124 4872 4204
rect 4872 4124 4952 4204
rect 4952 4124 5032 4204
rect 5032 4124 5112 4204
rect 32 158 112 238
rect 32 238 112 318
rect 32 318 112 398
rect 32 398 112 478
rect 32 478 112 558
rect 32 558 112 638
rect 32 638 112 718
rect 32 718 112 798
rect 32 798 112 878
rect 32 878 112 958
rect 32 958 112 1038
rect 32 1038 112 1118
rect 32 1118 112 1198
rect 32 1198 112 1278
rect 32 1278 112 1358
rect 32 1358 112 1438
rect 32 1438 112 1518
rect 32 1518 112 1598
rect 32 1598 112 1678
rect 32 1678 112 1758
rect 32 1758 112 1838
rect 32 1838 112 1918
rect 32 1918 112 1998
rect 32 1998 112 2078
rect 32 2078 112 2158
rect 32 2158 112 2238
rect 32 2238 112 2318
rect 32 2318 112 2398
rect 32 2398 112 2478
rect 32 2478 112 2558
rect 32 2558 112 2638
rect 32 2638 112 2718
rect 32 2718 112 2798
rect 32 2798 112 2878
rect 32 2878 112 2958
rect 32 2958 112 3038
rect 32 3038 112 3118
rect 32 3118 112 3198
rect 32 3198 112 3278
rect 32 3278 112 3358
rect 32 3358 112 3438
rect 32 3438 112 3518
rect 32 3518 112 3598
rect 32 3598 112 3678
rect 32 3678 112 3758
rect 32 3758 112 3838
rect 32 3838 112 3918
rect 32 3918 112 3998
rect 32 3998 112 4078
rect 5152 158 5232 238
rect 5152 238 5232 318
rect 5152 318 5232 398
rect 5152 398 5232 478
rect 5152 478 5232 558
rect 5152 558 5232 638
rect 5152 638 5232 718
rect 5152 718 5232 798
rect 5152 798 5232 878
rect 5152 878 5232 958
rect 5152 958 5232 1038
rect 5152 1038 5232 1118
rect 5152 1118 5232 1198
rect 5152 1198 5232 1278
rect 5152 1278 5232 1358
rect 5152 1358 5232 1438
rect 5152 1438 5232 1518
rect 5152 1518 5232 1598
rect 5152 1598 5232 1678
rect 5152 1678 5232 1758
rect 5152 1758 5232 1838
rect 5152 1838 5232 1918
rect 5152 1918 5232 1998
rect 5152 1998 5232 2078
rect 5152 2078 5232 2158
rect 5152 2158 5232 2238
rect 5152 2238 5232 2318
rect 5152 2318 5232 2398
rect 5152 2398 5232 2478
rect 5152 2478 5232 2558
rect 5152 2558 5232 2638
rect 5152 2638 5232 2718
rect 5152 2718 5232 2798
rect 5152 2798 5232 2878
rect 5152 2878 5232 2958
rect 5152 2958 5232 3038
rect 5152 3038 5232 3118
rect 5152 3118 5232 3198
rect 5152 3198 5232 3278
rect 5152 3278 5232 3358
rect 5152 3358 5232 3438
rect 5152 3438 5232 3518
rect 5152 3518 5232 3598
rect 5152 3598 5232 3678
rect 5152 3678 5232 3758
rect 5152 3758 5232 3838
rect 5152 3838 5232 3918
rect 5152 3918 5232 3998
rect 5152 3998 5232 4078
<< ptap >>
rect 0 0 5264 144
rect 0 4092 5264 4236
rect 0 0 144 4236
rect 5120 0 5264 4236
use SUNTR_RES8 XA1
transform 1 0 688 0 1 688
box 688 688 4576 3548
<< labels >>
flabel locali s 16 16 5248 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 4072 3438 4648 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
