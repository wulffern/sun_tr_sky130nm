magic
tech sky130B
magscale 1 2
timestamp 1669849200
<< checkpaint >>
rect 0 0 2520 1056
<< locali >>
rect 864 58 1032 118
rect 1032 58 1656 118
rect 1032 58 1092 118
rect 864 938 1032 998
rect 1032 938 1656 998
rect 1032 938 1092 998
rect 864 762 1032 822
rect 1032 762 1656 822
rect 1032 762 1092 822
rect 402 146 462 558
rect 432 850 600 910
rect 600 58 864 118
rect 600 58 660 910
rect 2088 146 2256 206
rect 2088 850 2256 910
rect 2256 146 2316 910
rect 834 234 894 470
rect 834 586 894 822
rect 1626 234 1686 470
rect 1626 586 1686 822
rect 1980 146 2196 206
rect 1548 762 1764 822
rect 756 938 972 998
<< poly >>
rect 324 158 2196 194
<< m3 >>
rect 1656 410 1836 486
rect 1836 498 2088 574
rect 1836 410 1912 574
rect 1548 0 1748 1056
rect 756 0 956 1056
rect 1548 0 1748 1056
rect 756 0 956 1056
use SUNTR_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTR_NCHDL MN2
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTR_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTR_PCHDL MP1_DMY
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTR_PCHDL MP2
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNTR_cut_M1M4_2x1 
transform 1 0 1548 0 1 410
box 1548 410 1748 486
use SUNTR_cut_M1M4_2x1 
transform 1 0 1980 0 1 498
box 1980 498 2180 574
use SUNTR_cut_M1M4_2x1 
transform 1 0 1548 0 1 234
box 1548 234 1748 310
use SUNTR_cut_M1M4_2x1 
transform 1 0 756 0 1 234
box 756 234 956 310
use SUNTR_cut_M1M4_2x1 
transform 1 0 756 0 1 410
box 756 410 956 486
<< labels >>
flabel locali s 1980 146 2196 206 0 FreeSans 400 0 0 0 C
port 1 nsew
flabel locali s 1548 762 1764 822 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 756 938 972 998 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel m3 s 1548 0 1748 1056 0 FreeSans 400 0 0 0 AVDD
port 4 nsew
flabel m3 s 756 0 956 1056 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
<< end >>
