magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 1260 3520
<< locali >>
rect 864 58 1032 118
rect 864 3402 1032 3462
rect 1032 58 1092 3462
rect 402 146 462 1966
rect 834 1642 894 1878
rect -108 132 108 220
rect 756 1642 972 1702
rect 324 146 540 206
rect 756 58 972 118
use SUNTR_NCHDLCM M0 
transform 1 0 0 0 1 0
box 0 0 1260 1760
use SUNTR_NCHDLCM M1 
transform 1 0 0 0 1 1760
box 0 1760 1260 3520
<< labels >>
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 756 1642 972 1702 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 756 58 972 118 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 3520
<< end >>
