* NGSPICE file created from SUNTR_PCHLA.ext - technology: sky130B

.subckt SUNTR_PCHLA D G S B
X0 D G S B sky130_fd_pr__pfet_01v8 ad=4.1472e+12p pd=2.496e+07u as=4.1472e+12p ps=2.496e+07u w=1.08e+06u l=360000u
X1 S G D B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X2 D G S B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X3 D G S B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X4 S G D B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X5 S G D B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X6 D G S B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
X7 S G D B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
C0 D S 0.82fF
C1 D G 0.53fF
C2 B S 0.76fF
C3 B G 2.44fF
C4 B D 0.52fF
C5 S 0 0.76fF
C6 G 0 0.54fF
C7 B 0 20.29fF
.ends
