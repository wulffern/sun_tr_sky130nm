magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 1260 4048
<< locali >>
rect 636 1642 864 1702
rect 636 3578 864 3638
rect 636 1642 696 3638
rect -108 132 108 220
rect 756 58 972 118
rect 756 3754 972 3814
rect 324 146 540 206
rect 324 3666 540 3726
rect 756 1642 972 1702
use SUNTR_NCHDLCM2 M0 
transform 1 0 0 0 1 0
box 0 0 1260 3520
use SUNTR_NCHDLA M1 
transform 1 0 0 0 1 3520
box 0 3520 1260 4048
<< labels >>
flabel locali s -108 132 108 220 0 FreeSans 400 0 0 0 B
port 6 nsew signal bidirectional
flabel locali s 756 58 972 118 0 FreeSans 400 0 0 0 S
port 4 nsew signal bidirectional
flabel locali s 756 3754 972 3814 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 324 3666 540 3726 0 FreeSans 400 0 0 0 CG
port 3 nsew signal bidirectional
flabel locali s 756 1642 972 1702 0 FreeSans 400 0 0 0 CS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 4048
<< end >>
