magic
tech sky130B
magscale 1 2
timestamp 1709161200
<< checkpaint >>
rect 0 0 1656 1056
<< m1 >>
rect 108 -44 1620 44
rect 1548 44 1620 132
rect 108 132 1476 220
rect 1548 132 1620 220
rect 108 220 180 308
rect 1548 220 1620 308
rect 108 308 180 396
rect 252 308 1620 396
rect 108 396 180 484
rect 1548 396 1620 484
rect 108 484 1476 572
rect 1548 484 1620 572
rect 108 572 180 660
rect 1548 572 1620 660
rect 108 660 180 748
rect 252 660 1620 748
rect 108 748 180 836
rect 108 836 1620 924
<< m2 >>
rect 108 -44 1620 44
rect 1548 44 1620 132
rect 108 132 1476 220
rect 1548 132 1620 220
rect 108 220 180 308
rect 1548 220 1620 308
rect 108 308 180 396
rect 252 308 1620 396
rect 108 396 180 484
rect 1548 396 1620 484
rect 108 484 1476 572
rect 1548 484 1620 572
rect 108 572 180 660
rect 1548 572 1620 660
rect 108 660 180 748
rect 252 660 1620 748
rect 108 748 180 836
rect 108 836 1620 924
<< locali >>
rect 108 -44 1620 44
rect 1548 44 1620 132
rect 108 132 1476 220
rect 1548 132 1620 220
rect 108 220 180 308
rect 1548 220 1620 308
rect 108 308 180 396
rect 252 308 1620 396
rect 108 396 180 484
rect 1548 396 1620 484
rect 108 484 1476 572
rect 1548 484 1620 572
rect 108 572 180 660
rect 1548 572 1620 660
rect 108 660 180 748
rect 252 660 1620 748
rect 108 748 180 836
rect 108 836 1620 924
<< v1 >>
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 1332 -35 1404 -26
rect 1332 -26 1404 -17
rect 1332 -17 1404 -8
rect 1332 -8 1404 0
rect 1332 0 1404 8
rect 1332 8 1404 17
rect 1332 17 1404 26
rect 1332 26 1404 35
rect 1404 -35 1476 -26
rect 1404 -26 1476 -17
rect 1404 -17 1476 -8
rect 1404 -8 1476 0
rect 1404 0 1476 8
rect 1404 8 1476 17
rect 1404 17 1476 26
rect 1404 26 1476 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 1332 316 1404 325
rect 1332 325 1404 334
rect 1332 334 1404 343
rect 1332 343 1404 352
rect 1332 352 1404 360
rect 1332 360 1404 369
rect 1332 369 1404 378
rect 1332 378 1404 387
rect 1404 316 1476 325
rect 1404 325 1476 334
rect 1404 334 1476 343
rect 1404 343 1476 352
rect 1404 352 1476 360
rect 1404 360 1476 369
rect 1404 369 1476 378
rect 1404 378 1476 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 1332 668 1404 677
rect 1332 677 1404 686
rect 1332 686 1404 695
rect 1332 695 1404 704
rect 1332 704 1404 712
rect 1332 712 1404 721
rect 1332 721 1404 730
rect 1332 730 1404 739
rect 1404 668 1476 677
rect 1404 677 1476 686
rect 1404 686 1476 695
rect 1404 695 1476 704
rect 1404 704 1476 712
rect 1404 712 1476 721
rect 1404 721 1476 730
rect 1404 730 1476 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 1332 -35 1404 -26
rect 1332 -26 1404 -17
rect 1332 -17 1404 -8
rect 1332 -8 1404 0
rect 1332 0 1404 8
rect 1332 8 1404 17
rect 1332 17 1404 26
rect 1332 26 1404 35
rect 1404 -35 1476 -26
rect 1404 -26 1476 -17
rect 1404 -17 1476 -8
rect 1404 -8 1476 0
rect 1404 0 1476 8
rect 1404 8 1476 17
rect 1404 17 1476 26
rect 1404 26 1476 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 1332 316 1404 325
rect 1332 325 1404 334
rect 1332 334 1404 343
rect 1332 343 1404 352
rect 1332 352 1404 360
rect 1332 360 1404 369
rect 1332 369 1404 378
rect 1332 378 1404 387
rect 1404 316 1476 325
rect 1404 325 1476 334
rect 1404 334 1476 343
rect 1404 343 1476 352
rect 1404 352 1476 360
rect 1404 360 1476 369
rect 1404 369 1476 378
rect 1404 378 1476 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 1332 668 1404 677
rect 1332 677 1404 686
rect 1332 686 1404 695
rect 1332 695 1404 704
rect 1332 704 1404 712
rect 1332 712 1404 721
rect 1332 721 1404 730
rect 1332 730 1404 739
rect 1404 668 1476 677
rect 1404 677 1476 686
rect 1404 686 1476 695
rect 1404 695 1476 704
rect 1404 704 1476 712
rect 1404 712 1476 721
rect 1404 721 1476 730
rect 1404 730 1476 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 1260 -35 1332 -26
rect 1260 -26 1332 -17
rect 1260 -17 1332 -8
rect 1260 -8 1332 0
rect 1260 0 1332 8
rect 1260 8 1332 17
rect 1260 17 1332 26
rect 1260 26 1332 35
rect 1332 -35 1404 -26
rect 1332 -26 1404 -17
rect 1332 -17 1404 -8
rect 1332 -8 1404 0
rect 1332 0 1404 8
rect 1332 8 1404 17
rect 1332 17 1404 26
rect 1332 26 1404 35
rect 1404 -35 1476 -26
rect 1404 -26 1476 -17
rect 1404 -17 1476 -8
rect 1404 -8 1476 0
rect 1404 0 1476 8
rect 1404 8 1476 17
rect 1404 17 1476 26
rect 1404 26 1476 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 1260 316 1332 325
rect 1260 325 1332 334
rect 1260 334 1332 343
rect 1260 343 1332 352
rect 1260 352 1332 360
rect 1260 360 1332 369
rect 1260 369 1332 378
rect 1260 378 1332 387
rect 1332 316 1404 325
rect 1332 325 1404 334
rect 1332 334 1404 343
rect 1332 343 1404 352
rect 1332 352 1404 360
rect 1332 360 1404 369
rect 1332 369 1404 378
rect 1332 378 1404 387
rect 1404 316 1476 325
rect 1404 325 1476 334
rect 1404 334 1476 343
rect 1404 343 1476 352
rect 1404 352 1476 360
rect 1404 360 1476 369
rect 1404 369 1476 378
rect 1404 378 1476 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 1260 668 1332 677
rect 1260 677 1332 686
rect 1260 686 1332 695
rect 1260 695 1332 704
rect 1260 704 1332 712
rect 1260 712 1332 721
rect 1260 721 1332 730
rect 1260 730 1332 739
rect 1332 668 1404 677
rect 1332 677 1404 686
rect 1332 686 1404 695
rect 1332 695 1404 704
rect 1332 704 1404 712
rect 1332 712 1404 721
rect 1332 721 1404 730
rect 1332 730 1404 739
rect 1404 668 1476 677
rect 1404 677 1476 686
rect 1404 686 1476 695
rect 1404 695 1476 704
rect 1404 704 1476 712
rect 1404 712 1476 721
rect 1404 721 1476 730
rect 1404 730 1476 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 1620 44
rect 108 -44 1620 44
rect 1548 44 1620 132
rect 108 132 1260 220
rect 1332 132 1476 220
rect 1548 132 1620 220
rect 108 220 180 308
rect 1548 220 1620 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 1620 396
rect 108 396 180 484
rect 1548 396 1620 484
rect 108 484 1476 572
rect 1548 484 1620 572
rect 108 572 180 660
rect 1548 572 1620 660
rect 108 660 180 748
rect 252 660 1620 748
rect 108 748 180 836
rect 108 836 1620 924
rect 108 836 1620 924
<< rm3 >>
rect 1260 132 1332 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 1620 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 836 1620 924 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1656 1056
<< end >>
