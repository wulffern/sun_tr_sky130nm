magic
tech sky130B
timestamp 1728046668
<< poly >>
rect 162 79 1098 97
<< locali >>
rect 378 117 828 147
rect 162 73 270 103
<< metal3 >>
rect 378 0 478 176
rect 774 0 874 176
use SUNTR_NCHDL  MN0
timestamp 1709161200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNTR_PCHDL  MP0
timestamp 1709161200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNTR_cut_M1M4_2x1  xcut0
timestamp 1709161200
transform 1 0 774 0 1 29
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut1
timestamp 1709161200
transform 1 0 378 0 1 29
box 0 0 100 38
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 200 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 117 486 147 0 FreeSans 200 0 0 0 Y
port 2 nsew signal bidirectional
flabel metal3 s 774 0 874 176 0 FreeSans 200 0 0 0 AVDD
port 3 nsew signal bidirectional
flabel metal3 s 378 0 478 176 0 FreeSans 200 0 0 0 AVSS
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
