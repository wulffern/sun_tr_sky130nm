magic
tech sky130B
magscale 1 2
timestamp 1672527600
<< checkpaint >>
rect 0 0 3536 4236
<< locali >>
rect 16 16 3520 128
rect 128 16 3408 128
rect 128 4108 3408 4220
rect 16 128 128 4108
rect 3408 128 3520 4108
rect 16 16 3520 128
rect 2344 3438 2920 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 168 32 248 112
rect 248 32 328 112
rect 328 32 408 112
rect 408 32 488 112
rect 488 32 568 112
rect 568 32 648 112
rect 648 32 728 112
rect 728 32 808 112
rect 808 32 888 112
rect 888 32 968 112
rect 968 32 1048 112
rect 1048 32 1128 112
rect 1128 32 1208 112
rect 1208 32 1288 112
rect 1288 32 1368 112
rect 1368 32 1448 112
rect 1448 32 1528 112
rect 1528 32 1608 112
rect 1608 32 1688 112
rect 1688 32 1768 112
rect 1768 32 1848 112
rect 1848 32 1928 112
rect 1928 32 2008 112
rect 2008 32 2088 112
rect 2088 32 2168 112
rect 2168 32 2248 112
rect 2248 32 2328 112
rect 2328 32 2408 112
rect 2408 32 2488 112
rect 2488 32 2568 112
rect 2568 32 2648 112
rect 2648 32 2728 112
rect 2728 32 2808 112
rect 2808 32 2888 112
rect 2888 32 2968 112
rect 2968 32 3048 112
rect 3048 32 3128 112
rect 3128 32 3208 112
rect 3208 32 3288 112
rect 3288 32 3368 112
rect 168 4124 248 4204
rect 248 4124 328 4204
rect 328 4124 408 4204
rect 408 4124 488 4204
rect 488 4124 568 4204
rect 568 4124 648 4204
rect 648 4124 728 4204
rect 728 4124 808 4204
rect 808 4124 888 4204
rect 888 4124 968 4204
rect 968 4124 1048 4204
rect 1048 4124 1128 4204
rect 1128 4124 1208 4204
rect 1208 4124 1288 4204
rect 1288 4124 1368 4204
rect 1368 4124 1448 4204
rect 1448 4124 1528 4204
rect 1528 4124 1608 4204
rect 1608 4124 1688 4204
rect 1688 4124 1768 4204
rect 1768 4124 1848 4204
rect 1848 4124 1928 4204
rect 1928 4124 2008 4204
rect 2008 4124 2088 4204
rect 2088 4124 2168 4204
rect 2168 4124 2248 4204
rect 2248 4124 2328 4204
rect 2328 4124 2408 4204
rect 2408 4124 2488 4204
rect 2488 4124 2568 4204
rect 2568 4124 2648 4204
rect 2648 4124 2728 4204
rect 2728 4124 2808 4204
rect 2808 4124 2888 4204
rect 2888 4124 2968 4204
rect 2968 4124 3048 4204
rect 3048 4124 3128 4204
rect 3128 4124 3208 4204
rect 3208 4124 3288 4204
rect 3288 4124 3368 4204
rect 32 158 112 238
rect 32 238 112 318
rect 32 318 112 398
rect 32 398 112 478
rect 32 478 112 558
rect 32 558 112 638
rect 32 638 112 718
rect 32 718 112 798
rect 32 798 112 878
rect 32 878 112 958
rect 32 958 112 1038
rect 32 1038 112 1118
rect 32 1118 112 1198
rect 32 1198 112 1278
rect 32 1278 112 1358
rect 32 1358 112 1438
rect 32 1438 112 1518
rect 32 1518 112 1598
rect 32 1598 112 1678
rect 32 1678 112 1758
rect 32 1758 112 1838
rect 32 1838 112 1918
rect 32 1918 112 1998
rect 32 1998 112 2078
rect 32 2078 112 2158
rect 32 2158 112 2238
rect 32 2238 112 2318
rect 32 2318 112 2398
rect 32 2398 112 2478
rect 32 2478 112 2558
rect 32 2558 112 2638
rect 32 2638 112 2718
rect 32 2718 112 2798
rect 32 2798 112 2878
rect 32 2878 112 2958
rect 32 2958 112 3038
rect 32 3038 112 3118
rect 32 3118 112 3198
rect 32 3198 112 3278
rect 32 3278 112 3358
rect 32 3358 112 3438
rect 32 3438 112 3518
rect 32 3518 112 3598
rect 32 3598 112 3678
rect 32 3678 112 3758
rect 32 3758 112 3838
rect 32 3838 112 3918
rect 32 3918 112 3998
rect 32 3998 112 4078
rect 3424 158 3504 238
rect 3424 238 3504 318
rect 3424 318 3504 398
rect 3424 398 3504 478
rect 3424 478 3504 558
rect 3424 558 3504 638
rect 3424 638 3504 718
rect 3424 718 3504 798
rect 3424 798 3504 878
rect 3424 878 3504 958
rect 3424 958 3504 1038
rect 3424 1038 3504 1118
rect 3424 1118 3504 1198
rect 3424 1198 3504 1278
rect 3424 1278 3504 1358
rect 3424 1358 3504 1438
rect 3424 1438 3504 1518
rect 3424 1518 3504 1598
rect 3424 1598 3504 1678
rect 3424 1678 3504 1758
rect 3424 1758 3504 1838
rect 3424 1838 3504 1918
rect 3424 1918 3504 1998
rect 3424 1998 3504 2078
rect 3424 2078 3504 2158
rect 3424 2158 3504 2238
rect 3424 2238 3504 2318
rect 3424 2318 3504 2398
rect 3424 2398 3504 2478
rect 3424 2478 3504 2558
rect 3424 2558 3504 2638
rect 3424 2638 3504 2718
rect 3424 2718 3504 2798
rect 3424 2798 3504 2878
rect 3424 2878 3504 2958
rect 3424 2958 3504 3038
rect 3424 3038 3504 3118
rect 3424 3118 3504 3198
rect 3424 3198 3504 3278
rect 3424 3278 3504 3358
rect 3424 3358 3504 3438
rect 3424 3438 3504 3518
rect 3424 3518 3504 3598
rect 3424 3598 3504 3678
rect 3424 3678 3504 3758
rect 3424 3758 3504 3838
rect 3424 3838 3504 3918
rect 3424 3918 3504 3998
rect 3424 3998 3504 4078
<< ptap >>
rect 0 0 3536 144
rect 0 4092 3536 4236
rect 0 0 144 4236
rect 3392 0 3536 4236
use SUNTR_RES4 XA1
transform 1 0 688 0 1 688
box 688 688 2848 3548
<< labels >>
flabel locali s 16 16 3520 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 2344 3438 2920 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
