magic
tech sky130A
magscale 1 2
timestamp 1711839600
<< checkpaint >>
rect 0 0 2520 352
<< locali >>
rect -108 146 540 206
rect 432 146 600 206
rect 600 58 864 118
rect 600 58 660 206
rect 432 146 600 206
rect 600 234 864 294
rect 600 146 660 294
rect 1656 58 1824 118
rect 1824 146 2088 206
rect 1824 58 1884 206
rect 1656 234 1824 294
rect 1824 146 2088 206
rect 1824 146 1884 294
rect 1980 146 2628 206
<< m3 >>
rect 1548 0 1748 352
rect 756 0 956 352
rect 1548 0 1748 352
rect 756 0 956 352
use SUNTR_NCHDL MN1 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_PCHDL MP1 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 234
box 1548 234 1748 310
use SUNTR_cut_M1M4_2x1 xcut1 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTR_cut_M1M4_2x1 xcut2 
transform 1 0 756 0 1 234
box 756 234 956 310
use SUNTR_cut_M1M4_2x1 xcut3 
transform 1 0 756 0 1 58
box 756 58 956 134
<< labels >>
flabel m3 s 1548 0 1748 352 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m3 s 756 0 956 352 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 352
<< end >>
