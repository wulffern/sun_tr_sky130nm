* NGSPICE file created from SUNTR_NCHLA.ext - technology: sky130B

.subckt SUNTR_NCHLA D G S B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=1.0368e+12p pd=6.24e+06u as=1.0368e+12p ps=6.24e+06u w=1.08e+06u l=360000u
X1 S G D B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=360000u
C0 M1/a_324_492# B 0.43fF $ **FLOATING
C1 S B 0.41fF
C2 G B 0.72fF
C3 M0/a_324_n36# B 0.43fF $ **FLOATING
.ends
