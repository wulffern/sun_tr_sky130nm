magic
tech sky130B
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 1296 2860
<< ppolyres >>
rect 360 -110 504 110
rect 792 -110 936 110
rect 360 110 504 330
rect 792 110 936 330
rect 360 330 504 550
rect 792 330 936 550
rect 360 550 504 770
rect 792 550 936 770
rect 360 770 504 990
rect 792 770 936 990
rect 360 990 504 1210
rect 792 990 936 1210
rect 360 1210 504 1430
rect 792 1210 936 1430
rect 360 1430 504 1650
rect 792 1430 936 1650
rect 360 1650 504 1870
rect 792 1650 936 1870
rect 360 1870 504 2090
rect 792 1870 936 2090
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
<< poly >>
rect -72 -110 72 110
rect 1224 -110 1368 110
rect -72 110 72 330
rect 1224 110 1368 330
rect -72 330 72 550
rect 1224 330 1368 550
rect -72 550 72 770
rect 1224 550 1368 770
rect -72 770 72 990
rect 1224 770 1368 990
rect -72 990 72 1210
rect 1224 990 1368 1210
rect -72 1210 72 1430
rect 1224 1210 1368 1430
rect -72 1430 72 1650
rect 1224 1430 1368 1650
rect -72 1650 72 1870
rect 1224 1650 1368 1870
rect -72 1870 72 2090
rect 1224 1870 1368 2090
rect -72 2090 72 2310
rect 1224 2090 1368 2310
rect -72 2310 72 2530
rect 1224 2310 1368 2530
<< xpolycontact >>
rect 360 -110 504 110
rect 792 -110 936 110
rect 360 110 504 330
rect 792 110 936 330
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
<< locali >>
rect 360 -110 936 110
rect 360 110 936 330
rect 360 2090 504 2310
rect 792 2090 936 2310
rect 360 2310 504 2530
rect 792 2310 936 2530
rect 360 2530 504 2750
rect 792 2530 936 2750
rect -72 2750 504 2970
rect -72 2750 504 2970
rect 792 2750 1368 2970
rect 792 2750 1368 2970
<< pwell >>
rect -72 -110 1368 2970
<< labels >>
flabel locali s -72 2750 504 2970 0 FreeSans 400 0 0 0 N
port 1 nsew
flabel locali s 792 2750 1368 2970 0 FreeSans 400 0 0 0 P
port 2 nsew
<< end >>
