magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 378 821 486 851
rect -54 66 54 110
rect 201 103 231 807
rect 162 73 270 103
rect 378 29 486 59
use SUNTR_NCHDL  M0
timestamp 1709161200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNTR_NCHDL  M1
timestamp 1709161200
transform 1 0 0 0 1 88
box -90 -66 630 242
use SUNTR_NCHDL  M2
timestamp 1709161200
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNTR_NCHDL  M3
timestamp 1709161200
transform 1 0 0 0 1 264
box -90 -66 630 242
use SUNTR_NCHDL  M4
timestamp 1709161200
transform 1 0 0 0 1 352
box -90 -66 630 242
use SUNTR_NCHDL  M5
timestamp 1709161200
transform 1 0 0 0 1 440
box -90 -66 630 242
use SUNTR_NCHDL  M6
timestamp 1709161200
transform 1 0 0 0 1 528
box -90 -66 630 242
use SUNTR_NCHDL  M7
timestamp 1709161200
transform 1 0 0 0 1 616
box -90 -66 630 242
use SUNTR_NCHDL  M8
timestamp 1709161200
transform 1 0 0 0 1 704
box -90 -66 630 242
<< labels >>
flabel locali s -54 66 54 110 0 FreeSans 200 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 378 821 486 851 0 FreeSans 200 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 73 270 103 0 FreeSans 200 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 378 29 486 59 0 FreeSans 200 0 0 0 S
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 630 880
<< end >>
