magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 2520 1056
<< locali >>
rect 834 586 894 822
rect 1626 234 1686 470
rect 864 410 1032 470
rect 1032 938 1656 998
rect 1032 410 1092 998
rect 204 850 432 910
rect 204 294 816 354
rect 204 294 264 910
rect 756 234 864 294
rect 864 234 1164 294
rect 1164 586 1656 646
rect 1164 234 1224 646
rect 324 146 540 206
rect 324 498 540 558
rect 756 410 972 470
<< poly >>
rect 324 158 2196 194
rect 324 510 2196 546
rect 324 862 2196 898
<< m3 >>
rect 1548 0 1748 1056
rect 756 0 956 1056
rect 1548 0 1748 1056
rect 756 0 956 1056
use SUNTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL MN2 
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTR_NCHDL MN1 
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTR_PCHDL MP1 
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTR_PCHDL MP0 
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTR_PCHDL MP2 
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNTR_cut_M1M4_2x1 xcut0 
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTR_cut_M1M4_2x1 xcut1 
transform 1 0 1548 0 1 762
box 1548 762 1748 838
use SUNTR_cut_M1M4_2x1 xcut2 
transform 1 0 756 0 1 58
box 756 58 956 134
use SUNTR_cut_M1M4_2x1 xcut3 
transform 1 0 756 0 1 938
box 756 938 956 1014
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 324 498 540 558 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 756 410 972 470 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel m3 s 1548 0 1748 1056 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 756 0 956 1056 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 1056
<< end >>
