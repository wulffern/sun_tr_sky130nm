magic
tech sky130B
magscale 1 2
timestamp 1709161200
<< checkpaint >>
rect 0 0 5400 1056
<< m1 >>
rect 108 -44 5364 44
rect 5292 44 5364 132
rect 108 132 5220 220
rect 5292 132 5364 220
rect 108 220 180 308
rect 5292 220 5364 308
rect 108 308 180 396
rect 252 308 5364 396
rect 108 396 180 484
rect 5292 396 5364 484
rect 108 484 5220 572
rect 5292 484 5364 572
rect 108 572 180 660
rect 5292 572 5364 660
rect 108 660 180 748
rect 252 660 5364 748
rect 108 748 180 836
rect 108 836 5364 924
<< m2 >>
rect 108 -44 5364 44
rect 5292 44 5364 132
rect 108 132 5220 220
rect 5292 132 5364 220
rect 108 220 180 308
rect 5292 220 5364 308
rect 108 308 180 396
rect 252 308 5364 396
rect 108 396 180 484
rect 5292 396 5364 484
rect 108 484 5220 572
rect 5292 484 5364 572
rect 108 572 180 660
rect 5292 572 5364 660
rect 108 660 180 748
rect 252 660 5364 748
rect 108 748 180 836
rect 108 836 5364 924
<< locali >>
rect 108 -44 5364 44
rect 5292 44 5364 132
rect 108 132 5220 220
rect 5292 132 5364 220
rect 108 220 180 308
rect 5292 220 5364 308
rect 108 308 180 396
rect 252 308 5364 396
rect 108 396 180 484
rect 5292 396 5364 484
rect 108 484 5220 572
rect 5292 484 5364 572
rect 108 572 180 660
rect 5292 572 5364 660
rect 108 660 180 748
rect 252 660 5364 748
rect 108 748 180 836
rect 108 836 5364 924
<< v1 >>
rect 5004 -35 5076 -26
rect 5004 -26 5076 -17
rect 5004 -17 5076 -8
rect 5004 -8 5076 0
rect 5004 0 5076 8
rect 5004 8 5076 17
rect 5004 17 5076 26
rect 5004 26 5076 35
rect 5076 -35 5148 -26
rect 5076 -26 5148 -17
rect 5076 -17 5148 -8
rect 5076 -8 5148 0
rect 5076 0 5148 8
rect 5076 8 5148 17
rect 5076 17 5148 26
rect 5076 26 5148 35
rect 5148 -35 5220 -26
rect 5148 -26 5220 -17
rect 5148 -17 5220 -8
rect 5148 -8 5220 0
rect 5148 0 5220 8
rect 5148 8 5220 17
rect 5148 17 5220 26
rect 5148 26 5220 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 5004 316 5076 325
rect 5004 325 5076 334
rect 5004 334 5076 343
rect 5004 343 5076 352
rect 5004 352 5076 360
rect 5004 360 5076 369
rect 5004 369 5076 378
rect 5004 378 5076 387
rect 5076 316 5148 325
rect 5076 325 5148 334
rect 5076 334 5148 343
rect 5076 343 5148 352
rect 5076 352 5148 360
rect 5076 360 5148 369
rect 5076 369 5148 378
rect 5076 378 5148 387
rect 5148 316 5220 325
rect 5148 325 5220 334
rect 5148 334 5220 343
rect 5148 343 5220 352
rect 5148 352 5220 360
rect 5148 360 5220 369
rect 5148 369 5220 378
rect 5148 378 5220 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 5004 668 5076 677
rect 5004 677 5076 686
rect 5004 686 5076 695
rect 5004 695 5076 704
rect 5004 704 5076 712
rect 5004 712 5076 721
rect 5004 721 5076 730
rect 5004 730 5076 739
rect 5076 668 5148 677
rect 5076 677 5148 686
rect 5076 686 5148 695
rect 5076 695 5148 704
rect 5076 704 5148 712
rect 5076 712 5148 721
rect 5076 721 5148 730
rect 5076 730 5148 739
rect 5148 668 5220 677
rect 5148 677 5220 686
rect 5148 686 5220 695
rect 5148 695 5220 704
rect 5148 704 5220 712
rect 5148 712 5220 721
rect 5148 721 5220 730
rect 5148 730 5220 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 5004 -35 5076 -26
rect 5004 -26 5076 -17
rect 5004 -17 5076 -8
rect 5004 -8 5076 0
rect 5004 0 5076 8
rect 5004 8 5076 17
rect 5004 17 5076 26
rect 5004 26 5076 35
rect 5076 -35 5148 -26
rect 5076 -26 5148 -17
rect 5076 -17 5148 -8
rect 5076 -8 5148 0
rect 5076 0 5148 8
rect 5076 8 5148 17
rect 5076 17 5148 26
rect 5076 26 5148 35
rect 5148 -35 5220 -26
rect 5148 -26 5220 -17
rect 5148 -17 5220 -8
rect 5148 -8 5220 0
rect 5148 0 5220 8
rect 5148 8 5220 17
rect 5148 17 5220 26
rect 5148 26 5220 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 5004 316 5076 325
rect 5004 325 5076 334
rect 5004 334 5076 343
rect 5004 343 5076 352
rect 5004 352 5076 360
rect 5004 360 5076 369
rect 5004 369 5076 378
rect 5004 378 5076 387
rect 5076 316 5148 325
rect 5076 325 5148 334
rect 5076 334 5148 343
rect 5076 343 5148 352
rect 5076 352 5148 360
rect 5076 360 5148 369
rect 5076 369 5148 378
rect 5076 378 5148 387
rect 5148 316 5220 325
rect 5148 325 5220 334
rect 5148 334 5220 343
rect 5148 343 5220 352
rect 5148 352 5220 360
rect 5148 360 5220 369
rect 5148 369 5220 378
rect 5148 378 5220 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 5004 668 5076 677
rect 5004 677 5076 686
rect 5004 686 5076 695
rect 5004 695 5076 704
rect 5004 704 5076 712
rect 5004 712 5076 721
rect 5004 721 5076 730
rect 5004 730 5076 739
rect 5076 668 5148 677
rect 5076 677 5148 686
rect 5076 686 5148 695
rect 5076 695 5148 704
rect 5076 704 5148 712
rect 5076 712 5148 721
rect 5076 721 5148 730
rect 5076 730 5148 739
rect 5148 668 5220 677
rect 5148 677 5220 686
rect 5148 686 5220 695
rect 5148 695 5220 704
rect 5148 704 5220 712
rect 5148 712 5220 721
rect 5148 721 5220 730
rect 5148 730 5220 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 5004 -35 5076 -26
rect 5004 -26 5076 -17
rect 5004 -17 5076 -8
rect 5004 -8 5076 0
rect 5004 0 5076 8
rect 5004 8 5076 17
rect 5004 17 5076 26
rect 5004 26 5076 35
rect 5076 -35 5148 -26
rect 5076 -26 5148 -17
rect 5076 -17 5148 -8
rect 5076 -8 5148 0
rect 5076 0 5148 8
rect 5076 8 5148 17
rect 5076 17 5148 26
rect 5076 26 5148 35
rect 5148 -35 5220 -26
rect 5148 -26 5220 -17
rect 5148 -17 5220 -8
rect 5148 -8 5220 0
rect 5148 0 5220 8
rect 5148 8 5220 17
rect 5148 17 5220 26
rect 5148 26 5220 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 5004 316 5076 325
rect 5004 325 5076 334
rect 5004 334 5076 343
rect 5004 343 5076 352
rect 5004 352 5076 360
rect 5004 360 5076 369
rect 5004 369 5076 378
rect 5004 378 5076 387
rect 5076 316 5148 325
rect 5076 325 5148 334
rect 5076 334 5148 343
rect 5076 343 5148 352
rect 5076 352 5148 360
rect 5076 360 5148 369
rect 5076 369 5148 378
rect 5076 378 5148 387
rect 5148 316 5220 325
rect 5148 325 5220 334
rect 5148 334 5220 343
rect 5148 343 5220 352
rect 5148 352 5220 360
rect 5148 360 5220 369
rect 5148 369 5220 378
rect 5148 378 5220 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 5004 668 5076 677
rect 5004 677 5076 686
rect 5004 686 5076 695
rect 5004 695 5076 704
rect 5004 704 5076 712
rect 5004 712 5076 721
rect 5004 721 5076 730
rect 5004 730 5076 739
rect 5076 668 5148 677
rect 5076 677 5148 686
rect 5076 686 5148 695
rect 5076 695 5148 704
rect 5076 704 5148 712
rect 5076 712 5148 721
rect 5076 721 5148 730
rect 5076 730 5148 739
rect 5148 668 5220 677
rect 5148 677 5220 686
rect 5148 686 5220 695
rect 5148 695 5220 704
rect 5148 704 5220 712
rect 5148 712 5220 721
rect 5148 721 5220 730
rect 5148 730 5220 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 5364 44
rect 108 -44 5364 44
rect 5292 44 5364 132
rect 108 132 5004 220
rect 5076 132 5220 220
rect 5292 132 5364 220
rect 108 220 180 308
rect 5292 220 5364 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 5364 396
rect 108 396 180 484
rect 5292 396 5364 484
rect 108 484 5220 572
rect 5292 484 5364 572
rect 108 572 180 660
rect 5292 572 5364 660
rect 108 660 180 748
rect 252 660 5364 748
rect 108 748 180 836
rect 108 836 5364 924
rect 108 836 5364 924
<< rm3 >>
rect 5004 132 5076 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 5364 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 836 5364 924 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5400 1056
<< end >>
