* NGSPICE file created from SUNTR_PCHDLCM2.ext - technology: sky130B

.subckt SUNTR_PCHDLCM2 D G S B
X0 M0/M7/S G S B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.2312e+12p ps=6.6e+06u w=1.08e+06u l=180000u
X1 D G M0/M7/S B sky130_fd_pr__pfet_01v8 ad=1.2312e+12p pd=6.6e+06u as=0p ps=0u w=1.08e+06u l=180000u
X2 M1/M7/S G D B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X3 S G M1/M7/S B sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
C0 B G 0.73fF
C1 B 0 6.00fF
.ends
