magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 144 205 252 235
rect 399 103 429 191
rect 360 73 468 103
rect 576 66 684 110
rect 144 29 252 59
use SUNTR_PCHDL  M0
timestamp 1709161200
transform 1 0 0 0 1 0
box 0 -66 720 242
use SUNTR_PCHDL  M7
timestamp 1709161200
transform 1 0 0 0 1 88
box 0 -66 720 242
<< labels >>
flabel locali s 576 66 684 110 0 FreeSans 200 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 144 205 252 235 0 FreeSans 200 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 360 73 468 103 0 FreeSans 200 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 144 29 252 59 0 FreeSans 200 0 0 0 S
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 630 264
<< end >>
