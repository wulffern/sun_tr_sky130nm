* NGSPICE file created from SUNTR_CNCHDLCM2.ext - technology: sky130B

.subckt SUNTR_CNCHDLCM2 D G CG S CS B
X0 M0/M0/M1/S G S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2312e+12p ps=6.6e+06u w=1.08e+06u l=180000u
X1 M0/M0/M2/S G M0/M0/M1/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X2 M0/M0/M3/S G M0/M0/M2/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X3 M0/M0/M4/S G M0/M0/M3/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X4 M0/M0/M5/S G M0/M0/M4/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X5 M0/M0/M6/S G M0/M0/M5/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X6 M0/M0/M7/S G M0/M0/M6/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X7 M0/M0/M8/S G M0/M0/M7/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X8 CS G M0/M0/M8/S B sky130_fd_pr__nfet_01v8 ad=2.4624e+12p pd=1.32e+07u as=0p ps=0u w=1.08e+06u l=180000u
X9 M0/M1/M1/S G CS B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X10 M0/M1/M2/S G M0/M1/M1/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X11 M0/M1/M3/S G M0/M1/M2/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X12 M0/M1/M4/S G M0/M1/M3/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X13 M0/M1/M5/S G M0/M1/M4/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X14 M0/M1/M6/S G M0/M1/M5/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X15 M0/M1/M7/S G M0/M1/M6/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X16 M0/M1/M8/S G M0/M1/M7/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X17 S G M0/M1/M8/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X18 D CG CS B sky130_fd_pr__nfet_01v8 ad=7.56025e+11p pd=3.565e+06u as=0p ps=0u w=1.08e+06u l=180000u
X19 CS CG D B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
C0 CG B 0.47fF
C1 G B 4.10fF
C2 CS B 0.51fF
C3 S B 1.16fF
.ends
