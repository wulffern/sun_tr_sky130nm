* NGSPICE file created from SUNTR_NCHDLCM.ext - technology: sky130B

.subckt SUNTR_NCHDLCM D G S B
X0 M1/S G S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.156e+11p ps=3.3e+06u w=1.08e+06u l=180000u
X1 M2/S G M1/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X2 M3/S G M2/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X3 M5/S G M4/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X4 M4/S G M3/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X5 M6/S G M5/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X6 M7/S G M6/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X7 M8/S G M7/S B sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.08e+06u l=180000u
X8 D G M8/S B sky130_fd_pr__nfet_01v8 ad=6.156e+11p pd=3.3e+06u as=0p ps=0u w=1.08e+06u l=180000u
C0 G B 2.15fF
.ends
