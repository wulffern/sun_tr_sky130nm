magic
tech sky130B
timestamp 1728046668
<< poly >>
rect 162 255 1098 273
rect 162 79 1098 97
<< locali >>
rect 378 469 828 499
rect 162 425 270 455
rect 990 425 1098 455
rect 417 323 447 411
rect 813 323 843 411
rect 378 293 882 323
rect 162 249 270 279
rect 417 117 447 235
rect 162 73 270 103
rect 714 59 744 293
rect 714 29 828 59
<< metal3 >>
rect 378 0 478 528
rect 774 0 874 528
use SUNTR_NCHDL  MN0
timestamp 1709161200
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNTR_NCHDL  MN1
timestamp 1709161200
transform 1 0 0 0 1 352
box -90 -66 630 242
use SUNTR_NCHDL  MN2
timestamp 1709161200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNTR_PCHDL  MP0
timestamp 1709161200
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNTR_PCHDL  MP1
timestamp 1709161200
transform 1 0 630 0 1 352
box 0 -66 720 242
use SUNTR_PCHDL  MP2
timestamp 1709161200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNTR_cut_M1M4_2x1  xcut0
timestamp 1709161200
transform 1 0 774 0 1 117
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut1
timestamp 1709161200
transform 1 0 774 0 1 205
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut2
timestamp 1709161200
transform 1 0 378 0 1 29
box 0 0 100 38
<< labels >>
flabel locali s 162 249 270 279 0 FreeSans 200 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 990 425 1098 455 0 FreeSans 200 0 0 0 CN
port 3 nsew signal bidirectional
flabel locali s 162 425 270 455 0 FreeSans 200 0 0 0 C
port 2 nsew signal bidirectional
flabel locali s 162 73 270 103 0 FreeSans 200 0 0 0 RN
port 4 nsew signal bidirectional
flabel locali s 378 469 486 499 0 FreeSans 200 0 0 0 Y
port 5 nsew signal bidirectional
flabel metal3 s 774 0 874 528 0 FreeSans 200 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel metal3 s 378 0 478 528 0 FreeSans 200 0 0 0 AVSS
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 528
<< end >>
