magic
tech sky130A
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect -1440 -1440 16560 7072
<< locali >>
rect 15640 -720 15840 6352
rect -720 -720 15840 -520
rect -720 6152 15840 6352
rect -720 -720 -520 6352
rect 15640 -720 15840 6352
rect 16360 -1440 16560 7072
rect -1440 -1440 16560 -1240
rect -1440 6872 16560 7072
rect -1440 -1440 -1240 7072
rect 16360 -1440 16560 7072
<< m3 >>
rect 756 -720 956 352
rect 756 -720 956 704
rect 756 -720 956 1056
rect 4084 -720 4284 352
rect 4084 -720 4284 704
rect 4084 -720 4284 1408
rect 4084 -720 4284 2816
rect 4084 -720 4284 5632
rect 5796 -720 5996 352
rect 5796 -720 5996 1056
rect 9124 -720 9324 352
rect 9124 -720 9324 1056
rect 9124 -720 9324 1760
rect 9124 -720 9324 2816
rect 9124 -720 9324 3872
rect 10836 -720 11036 352
rect 10836 -720 11036 2112
rect 14164 -720 14364 352
rect 14164 -720 14364 1056
rect 14164 -720 14364 2464
rect 14164 -720 14364 3520
rect 1548 -1440 1748 352
rect 1548 -1440 1748 704
rect 1548 -1440 1748 1056
rect 3292 -1440 3492 352
rect 3292 -1440 3492 704
rect 3292 -1440 3492 1408
rect 3292 -1440 3492 2816
rect 3292 -1440 3492 5632
rect 6588 -1440 6788 352
rect 6588 -1440 6788 1056
rect 8332 -1440 8532 352
rect 8332 -1440 8532 1056
rect 8332 -1440 8532 1760
rect 8332 -1440 8532 2816
rect 8332 -1440 8532 3872
rect 11628 -1440 11828 352
rect 11628 -1440 11828 2112
rect 13372 -1440 13572 352
rect 13372 -1440 13572 3520
use SUNTR_TAPCELLB_CV XA0
transform 1 0 0 0 1 0
box 0 0 2520 352
use SUNTR_TIEH_CV XA1
transform 1 0 0 0 1 352
box 0 352 2520 704
use SUNTR_TIEL_CV XA2
transform 1 0 0 0 1 704
box 0 704 2520 1056
use SUNTR_TAPCELLB_CV XB0
transform -1 0 5040 0 1 0
box 5040 0 7560 352
use SUNTR_IVX1_CV XB3
transform -1 0 5040 0 1 352
box 5040 352 7560 704
use SUNTR_IVX2_CV XB4
transform -1 0 5040 0 1 704
box 5040 704 7560 1408
use SUNTR_IVX4_CV XB5
transform -1 0 5040 0 1 1408
box 5040 1408 7560 2816
use SUNTR_IVX8_CV XB6
transform -1 0 5040 0 1 2816
box 5040 2816 7560 5632
use SUNTR_TAPCELLB_CV XC0
transform 1 0 5040 0 1 0
box 5040 0 7560 352
use SUNTR_BFX1_CV XC7
transform 1 0 5040 0 1 352
box 5040 352 7560 1056
use SUNTR_TAPCELLB_CV XD0
transform -1 0 10080 0 1 0
box 10080 0 12600 352
use SUNTR_NRX1_CV XD8
transform -1 0 10080 0 1 352
box 10080 352 12600 1056
use SUNTR_NDX1_CV XD9
transform -1 0 10080 0 1 1056
box 10080 1056 12600 1760
use SUNTR_ORX1_CV XD10
transform -1 0 10080 0 1 1760
box 10080 1760 12600 2816
use SUNTR_ANX1_CV XD11
transform -1 0 10080 0 1 2816
box 10080 2816 12600 3872
use SUNTR_TAPCELLB_CV XE0
transform 1 0 10080 0 1 0
box 10080 0 12600 352
use SUNTR_SCX1_CV XE12
transform 1 0 10080 0 1 352
box 10080 352 12600 2112
use SUNTR_TAPCELLB_CV XF0
transform -1 0 15120 0 1 0
box 15120 0 17640 352
use SUNTR_SWX2_CV XF13
transform -1 0 15120 0 1 352
box 15120 352 17640 1056
use SUNTR_SWX4_CV XF14
transform -1 0 15120 0 1 1056
box 15120 1056 17640 2464
use SUNTR_TGPD_CV XF15
transform -1 0 15120 0 1 2464
box 15120 2464 17640 3520
use SUNTR_cut_M1M4_2x2 
transform 1 0 756 0 1 -720
box 756 -720 956 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 756 0 1 -720
box 756 -720 956 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 756 0 1 -720
box 756 -720 956 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 4084 0 1 -720
box 4084 -720 4284 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 5796 0 1 -720
box 5796 -720 5996 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 5796 0 1 -720
box 5796 -720 5996 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 9124 0 1 -720
box 9124 -720 9324 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 10836 0 1 -720
box 10836 -720 11036 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 10836 0 1 -720
box 10836 -720 11036 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 14164 0 1 -720
box 14164 -720 14364 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 14164 0 1 -720
box 14164 -720 14364 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 14164 0 1 -720
box 14164 -720 14364 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 14164 0 1 -720
box 14164 -720 14364 -520
use SUNTR_cut_M1M4_2x2 
transform 1 0 1548 0 1 -1440
box 1548 -1440 1748 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 1548 0 1 -1440
box 1548 -1440 1748 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 1548 0 1 -1440
box 1548 -1440 1748 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 3292 0 1 -1440
box 3292 -1440 3492 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 6588 0 1 -1440
box 6588 -1440 6788 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 6588 0 1 -1440
box 6588 -1440 6788 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 8332 0 1 -1440
box 8332 -1440 8532 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 11628 0 1 -1440
box 11628 -1440 11828 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 11628 0 1 -1440
box 11628 -1440 11828 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 13372 0 1 -1440
box 13372 -1440 13572 -1240
use SUNTR_cut_M1M4_2x2 
transform 1 0 13372 0 1 -1440
box 13372 -1440 13572 -1240
<< labels >>
flabel locali s 15640 -720 15840 6352 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 16360 -1440 16560 7072 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
<< end >>
