magic
tech sky130A
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 8720 4236
<< locali >>
rect 16 16 8704 128
rect 16 16 8704 128
rect 16 16 128 4220
rect 16 4108 8704 4220
rect 8592 16 8704 4220
rect 16 16 8704 128
rect 7528 3438 8104 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 40 32 120 112
rect 120 32 200 112
rect 200 32 280 112
rect 280 32 360 112
rect 360 32 440 112
rect 440 32 520 112
rect 520 32 600 112
rect 600 32 680 112
rect 680 32 760 112
rect 760 32 840 112
rect 840 32 920 112
rect 920 32 1000 112
rect 1000 32 1080 112
rect 1080 32 1160 112
rect 1160 32 1240 112
rect 1240 32 1320 112
rect 1320 32 1400 112
rect 1400 32 1480 112
rect 1480 32 1560 112
rect 1560 32 1640 112
rect 1640 32 1720 112
rect 1720 32 1800 112
rect 1800 32 1880 112
rect 1880 32 1960 112
rect 1960 32 2040 112
rect 2040 32 2120 112
rect 2120 32 2200 112
rect 2200 32 2280 112
rect 2280 32 2360 112
rect 2360 32 2440 112
rect 2440 32 2520 112
rect 2520 32 2600 112
rect 2600 32 2680 112
rect 2680 32 2760 112
rect 2760 32 2840 112
rect 2840 32 2920 112
rect 2920 32 3000 112
rect 3000 32 3080 112
rect 3080 32 3160 112
rect 3160 32 3240 112
rect 3240 32 3320 112
rect 3320 32 3400 112
rect 3400 32 3480 112
rect 3480 32 3560 112
rect 3560 32 3640 112
rect 3640 32 3720 112
rect 3720 32 3800 112
rect 3800 32 3880 112
rect 3880 32 3960 112
rect 3960 32 4040 112
rect 4040 32 4120 112
rect 4120 32 4200 112
rect 4200 32 4280 112
rect 4280 32 4360 112
rect 4360 32 4440 112
rect 4440 32 4520 112
rect 4520 32 4600 112
rect 4600 32 4680 112
rect 4680 32 4760 112
rect 4760 32 4840 112
rect 4840 32 4920 112
rect 4920 32 5000 112
rect 5000 32 5080 112
rect 5080 32 5160 112
rect 5160 32 5240 112
rect 5240 32 5320 112
rect 5320 32 5400 112
rect 5400 32 5480 112
rect 5480 32 5560 112
rect 5560 32 5640 112
rect 5640 32 5720 112
rect 5720 32 5800 112
rect 5800 32 5880 112
rect 5880 32 5960 112
rect 5960 32 6040 112
rect 6040 32 6120 112
rect 6120 32 6200 112
rect 6200 32 6280 112
rect 6280 32 6360 112
rect 6360 32 6440 112
rect 6440 32 6520 112
rect 6520 32 6600 112
rect 6600 32 6680 112
rect 6680 32 6760 112
rect 6760 32 6840 112
rect 6840 32 6920 112
rect 6920 32 7000 112
rect 7000 32 7080 112
rect 7080 32 7160 112
rect 7160 32 7240 112
rect 7240 32 7320 112
rect 7320 32 7400 112
rect 7400 32 7480 112
rect 7480 32 7560 112
rect 7560 32 7640 112
rect 7640 32 7720 112
rect 7720 32 7800 112
rect 7800 32 7880 112
rect 7880 32 7960 112
rect 7960 32 8040 112
rect 8040 32 8120 112
rect 8120 32 8200 112
rect 8200 32 8280 112
rect 8280 32 8360 112
rect 8360 32 8440 112
rect 8440 32 8520 112
rect 8520 32 8600 112
rect 8600 32 8680 112
rect 32 38 112 118
rect 32 118 112 198
rect 32 198 112 278
rect 32 278 112 358
rect 32 358 112 438
rect 32 438 112 518
rect 32 518 112 598
rect 32 598 112 678
rect 32 678 112 758
rect 32 758 112 838
rect 32 838 112 918
rect 32 918 112 998
rect 32 998 112 1078
rect 32 1078 112 1158
rect 32 1158 112 1238
rect 32 1238 112 1318
rect 32 1318 112 1398
rect 32 1398 112 1478
rect 32 1478 112 1558
rect 32 1558 112 1638
rect 32 1638 112 1718
rect 32 1718 112 1798
rect 32 1798 112 1878
rect 32 1878 112 1958
rect 32 1958 112 2038
rect 32 2038 112 2118
rect 32 2118 112 2198
rect 32 2198 112 2278
rect 32 2278 112 2358
rect 32 2358 112 2438
rect 32 2438 112 2518
rect 32 2518 112 2598
rect 32 2598 112 2678
rect 32 2678 112 2758
rect 32 2758 112 2838
rect 32 2838 112 2918
rect 32 2918 112 2998
rect 32 2998 112 3078
rect 32 3078 112 3158
rect 32 3158 112 3238
rect 32 3238 112 3318
rect 32 3318 112 3398
rect 32 3398 112 3478
rect 32 3478 112 3558
rect 32 3558 112 3638
rect 32 3638 112 3718
rect 32 3718 112 3798
rect 32 3798 112 3878
rect 32 3878 112 3958
rect 32 3958 112 4038
rect 32 4038 112 4118
rect 32 4118 112 4198
rect 40 4124 120 4204
rect 120 4124 200 4204
rect 200 4124 280 4204
rect 280 4124 360 4204
rect 360 4124 440 4204
rect 440 4124 520 4204
rect 520 4124 600 4204
rect 600 4124 680 4204
rect 680 4124 760 4204
rect 760 4124 840 4204
rect 840 4124 920 4204
rect 920 4124 1000 4204
rect 1000 4124 1080 4204
rect 1080 4124 1160 4204
rect 1160 4124 1240 4204
rect 1240 4124 1320 4204
rect 1320 4124 1400 4204
rect 1400 4124 1480 4204
rect 1480 4124 1560 4204
rect 1560 4124 1640 4204
rect 1640 4124 1720 4204
rect 1720 4124 1800 4204
rect 1800 4124 1880 4204
rect 1880 4124 1960 4204
rect 1960 4124 2040 4204
rect 2040 4124 2120 4204
rect 2120 4124 2200 4204
rect 2200 4124 2280 4204
rect 2280 4124 2360 4204
rect 2360 4124 2440 4204
rect 2440 4124 2520 4204
rect 2520 4124 2600 4204
rect 2600 4124 2680 4204
rect 2680 4124 2760 4204
rect 2760 4124 2840 4204
rect 2840 4124 2920 4204
rect 2920 4124 3000 4204
rect 3000 4124 3080 4204
rect 3080 4124 3160 4204
rect 3160 4124 3240 4204
rect 3240 4124 3320 4204
rect 3320 4124 3400 4204
rect 3400 4124 3480 4204
rect 3480 4124 3560 4204
rect 3560 4124 3640 4204
rect 3640 4124 3720 4204
rect 3720 4124 3800 4204
rect 3800 4124 3880 4204
rect 3880 4124 3960 4204
rect 3960 4124 4040 4204
rect 4040 4124 4120 4204
rect 4120 4124 4200 4204
rect 4200 4124 4280 4204
rect 4280 4124 4360 4204
rect 4360 4124 4440 4204
rect 4440 4124 4520 4204
rect 4520 4124 4600 4204
rect 4600 4124 4680 4204
rect 4680 4124 4760 4204
rect 4760 4124 4840 4204
rect 4840 4124 4920 4204
rect 4920 4124 5000 4204
rect 5000 4124 5080 4204
rect 5080 4124 5160 4204
rect 5160 4124 5240 4204
rect 5240 4124 5320 4204
rect 5320 4124 5400 4204
rect 5400 4124 5480 4204
rect 5480 4124 5560 4204
rect 5560 4124 5640 4204
rect 5640 4124 5720 4204
rect 5720 4124 5800 4204
rect 5800 4124 5880 4204
rect 5880 4124 5960 4204
rect 5960 4124 6040 4204
rect 6040 4124 6120 4204
rect 6120 4124 6200 4204
rect 6200 4124 6280 4204
rect 6280 4124 6360 4204
rect 6360 4124 6440 4204
rect 6440 4124 6520 4204
rect 6520 4124 6600 4204
rect 6600 4124 6680 4204
rect 6680 4124 6760 4204
rect 6760 4124 6840 4204
rect 6840 4124 6920 4204
rect 6920 4124 7000 4204
rect 7000 4124 7080 4204
rect 7080 4124 7160 4204
rect 7160 4124 7240 4204
rect 7240 4124 7320 4204
rect 7320 4124 7400 4204
rect 7400 4124 7480 4204
rect 7480 4124 7560 4204
rect 7560 4124 7640 4204
rect 7640 4124 7720 4204
rect 7720 4124 7800 4204
rect 7800 4124 7880 4204
rect 7880 4124 7960 4204
rect 7960 4124 8040 4204
rect 8040 4124 8120 4204
rect 8120 4124 8200 4204
rect 8200 4124 8280 4204
rect 8280 4124 8360 4204
rect 8360 4124 8440 4204
rect 8440 4124 8520 4204
rect 8520 4124 8600 4204
rect 8600 4124 8680 4204
rect 8608 38 8688 118
rect 8608 118 8688 198
rect 8608 198 8688 278
rect 8608 278 8688 358
rect 8608 358 8688 438
rect 8608 438 8688 518
rect 8608 518 8688 598
rect 8608 598 8688 678
rect 8608 678 8688 758
rect 8608 758 8688 838
rect 8608 838 8688 918
rect 8608 918 8688 998
rect 8608 998 8688 1078
rect 8608 1078 8688 1158
rect 8608 1158 8688 1238
rect 8608 1238 8688 1318
rect 8608 1318 8688 1398
rect 8608 1398 8688 1478
rect 8608 1478 8688 1558
rect 8608 1558 8688 1638
rect 8608 1638 8688 1718
rect 8608 1718 8688 1798
rect 8608 1798 8688 1878
rect 8608 1878 8688 1958
rect 8608 1958 8688 2038
rect 8608 2038 8688 2118
rect 8608 2118 8688 2198
rect 8608 2198 8688 2278
rect 8608 2278 8688 2358
rect 8608 2358 8688 2438
rect 8608 2438 8688 2518
rect 8608 2518 8688 2598
rect 8608 2598 8688 2678
rect 8608 2678 8688 2758
rect 8608 2758 8688 2838
rect 8608 2838 8688 2918
rect 8608 2918 8688 2998
rect 8608 2998 8688 3078
rect 8608 3078 8688 3158
rect 8608 3158 8688 3238
rect 8608 3238 8688 3318
rect 8608 3318 8688 3398
rect 8608 3398 8688 3478
rect 8608 3478 8688 3558
rect 8608 3558 8688 3638
rect 8608 3638 8688 3718
rect 8608 3718 8688 3798
rect 8608 3798 8688 3878
rect 8608 3878 8688 3958
rect 8608 3958 8688 4038
rect 8608 4038 8688 4118
rect 8608 4118 8688 4198
<< ptap >>
rect 0 0 8720 144
rect 0 0 144 4236
rect 0 4092 8720 4236
rect 8576 0 8720 4236
use SUNTR_RES16 XA1
transform 1 0 688 0 1 688
box 688 688 8032 3548
<< labels >>
flabel locali s 16 16 8704 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 7528 3438 8104 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
