magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 378 2581 486 2611
rect 216 2537 330 2567
rect 300 2435 330 2537
rect 300 2405 486 2435
rect 912 2361 1044 2391
rect 162 2009 270 2039
rect 216 1833 270 1863
rect 240 1803 330 1833
rect 300 1335 330 1803
rect 432 1349 546 1379
rect 216 1305 330 1335
rect 300 675 330 1305
rect 516 1027 546 1349
rect 432 997 546 1027
rect 912 983 942 2361
rect 912 953 1044 983
rect 912 675 942 953
rect 990 777 1098 807
rect 300 645 432 675
rect 828 645 942 675
rect 990 601 1044 631
rect 912 571 1020 601
rect 912 323 942 571
rect 828 293 942 323
rect 162 249 270 279
<< metal1 >>
rect 828 2581 942 2611
rect 432 2405 546 2435
rect 102 2009 216 2039
rect 102 455 132 2009
rect 516 1907 546 2405
rect 912 2215 942 2581
rect 912 2185 1044 2215
rect 432 1877 546 1907
rect 1044 1833 1158 1863
rect 912 1657 1044 1687
rect 912 1555 942 1657
rect 828 1525 942 1555
rect 216 1481 330 1511
rect 300 1379 330 1481
rect 300 1349 432 1379
rect 912 1159 942 1525
rect 1128 1335 1158 1833
rect 1044 1305 1158 1335
rect 912 1129 1044 1159
rect 216 953 270 983
rect 240 923 330 953
rect 300 499 330 923
rect 300 469 432 499
rect 102 425 216 455
rect 1128 323 1158 1305
rect 828 293 1158 323
<< metal2 >>
rect 216 2361 340 2399
rect 302 1871 340 2361
rect 302 1833 1044 1871
<< metal3 >>
rect 378 0 478 2640
rect 774 0 874 2640
use SUNTR_TAPCELLB_CV  XA0
timestamp 1728046668
transform 1 0 0 0 1 0
box -90 -66 1350 242
use SUNTR_NDX1_CV  XA1
timestamp 1728046668
transform 1 0 0 0 1 176
box -90 -66 1350 418
use SUNTR_IVX1_CV  XA2
timestamp 1728046668
transform 1 0 0 0 1 528
box -90 -66 1350 242
use SUNTR_IVTRIX1_CV  XA3
timestamp 1728046668
transform 1 0 0 0 1 704
box -90 -66 1350 418
use SUNTR_IVTRIX1_CV  XA4
timestamp 1728046668
transform 1 0 0 0 1 1056
box -90 -66 1350 418
use SUNTR_IVX1_CV  XA5
timestamp 1728046668
transform 1 0 0 0 1 1408
box -90 -66 1350 242
use SUNTR_IVTRIX1_CV  XA6
timestamp 1728046668
transform 1 0 0 0 1 1584
box -90 -66 1350 418
use SUNTR_NDTRIX1_CV  XA7
timestamp 1728046668
transform 1 0 0 0 1 1936
box -90 -66 1350 594
use SUNTR_IVX1_CV  XA8
timestamp 1728046668
transform 1 0 0 0 1 2464
box -90 -66 1350 242
use SUNTR_cut_M1M2_2x1  xcut0
timestamp 1709161200
transform 1 0 990 0 1 1305
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut1
timestamp 1709161200
transform 1 0 990 0 1 1833
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut2
timestamp 1709161200
transform 1 0 774 0 1 293
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut3
timestamp 1709161200
transform 1 0 162 0 1 953
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut4
timestamp 1709161200
transform 1 0 378 0 1 469
box 0 0 92 34
use SUNTR_cut_M1M3_2x1  xcut5
timestamp 1709161200
transform 1 0 162 0 1 2361
box 0 0 100 38
use SUNTR_cut_M1M3_2x1  xcut6
timestamp 1709161200
transform 1 0 990 0 1 1833
box 0 0 100 38
use SUNTR_cut_M1M2_2x1  xcut7
timestamp 1709161200
transform 1 0 378 0 1 1877
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut8
timestamp 1709161200
transform 1 0 378 0 1 2405
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut9
timestamp 1709161200
transform 1 0 162 0 1 1481
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut10
timestamp 1709161200
transform 1 0 378 0 1 1349
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut11
timestamp 1709161200
transform 1 0 774 0 1 1525
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut12
timestamp 1709161200
transform 1 0 990 0 1 1129
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut13
timestamp 1709161200
transform 1 0 990 0 1 1657
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut14
timestamp 1709161200
transform 1 0 774 0 1 2581
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut15
timestamp 1709161200
transform 1 0 990 0 1 2185
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut16
timestamp 1709161200
transform 1 0 162 0 1 425
box 0 0 92 34
use SUNTR_cut_M1M2_2x1  xcut17
timestamp 1709161200
transform 1 0 162 0 1 2009
box 0 0 92 34
<< labels >>
flabel locali s 990 777 1098 807 0 FreeSans 200 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 249 270 279 0 FreeSans 200 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 2581 486 2611 0 FreeSans 200 0 0 0 Q
port 4 nsew signal bidirectional
flabel locali s 378 2405 486 2435 0 FreeSans 200 0 0 0 QN
port 5 nsew signal bidirectional
flabel metal3 s 774 0 874 2640 0 FreeSans 200 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel metal3 s 378 0 478 2640 0 FreeSans 200 0 0 0 AVSS
port 7 nsew signal bidirectional
flabel locali s 162 2009 270 2039 0 FreeSans 200 0 0 0 RN
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 2640
<< end >>
