magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 300 117 432 147
rect 828 117 942 147
rect 300 103 330 117
rect -54 73 330 103
rect 300 59 330 73
rect 912 103 942 117
rect 912 73 1314 103
rect 912 59 942 73
rect 300 29 432 59
rect 828 29 942 59
<< metal3 >>
rect 378 0 478 176
rect 774 0 874 176
use SUNTR_NCHDL  MN1
timestamp 1709161200
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNTR_PCHDL  MP1
timestamp 1709161200
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNTR_cut_M1M4_2x1  xcut0
timestamp 1709161200
transform 1 0 774 0 1 117
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut1
timestamp 1709161200
transform 1 0 774 0 1 29
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut2
timestamp 1709161200
transform 1 0 378 0 1 117
box 0 0 100 38
use SUNTR_cut_M1M4_2x1  xcut3
timestamp 1709161200
transform 1 0 378 0 1 29
box 0 0 100 38
<< labels >>
flabel metal3 s 774 0 874 176 0 FreeSans 200 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal3 s 378 0 478 176 0 FreeSans 200 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
