magic
tech sky130A
magscale 1 2
timestamp 1711839600
<< checkpaint >>
rect 0 0 2952 1056
<< m1 >>
rect 108 -44 2916 44
rect 2844 44 2916 132
rect 108 132 2772 220
rect 2844 132 2916 220
rect 108 220 180 308
rect 2844 220 2916 308
rect 108 308 180 396
rect 252 308 2916 396
rect 108 396 180 484
rect 2844 396 2916 484
rect 108 484 2772 572
rect 2844 484 2916 572
rect 108 572 180 660
rect 2844 572 2916 660
rect 108 660 180 748
rect 252 660 2916 748
rect 108 748 180 836
rect 108 836 2916 924
<< m2 >>
rect 108 -44 2916 44
rect 2844 44 2916 132
rect 108 132 2772 220
rect 2844 132 2916 220
rect 108 220 180 308
rect 2844 220 2916 308
rect 108 308 180 396
rect 252 308 2916 396
rect 108 396 180 484
rect 2844 396 2916 484
rect 108 484 2772 572
rect 2844 484 2916 572
rect 108 572 180 660
rect 2844 572 2916 660
rect 108 660 180 748
rect 252 660 2916 748
rect 108 748 180 836
rect 108 836 2916 924
<< locali >>
rect 108 -44 2916 44
rect 2844 44 2916 132
rect 108 132 2772 220
rect 2844 132 2916 220
rect 108 220 180 308
rect 2844 220 2916 308
rect 108 308 180 396
rect 252 308 2916 396
rect 108 396 180 484
rect 2844 396 2916 484
rect 108 484 2772 572
rect 2844 484 2916 572
rect 108 572 180 660
rect 2844 572 2916 660
rect 108 660 180 748
rect 252 660 2916 748
rect 108 748 180 836
rect 108 836 2916 924
<< v1 >>
rect 2556 -35 2628 -26
rect 2556 -26 2628 -17
rect 2556 -17 2628 -8
rect 2556 -8 2628 0
rect 2556 0 2628 8
rect 2556 8 2628 17
rect 2556 17 2628 26
rect 2556 26 2628 35
rect 2628 -35 2700 -26
rect 2628 -26 2700 -17
rect 2628 -17 2700 -8
rect 2628 -8 2700 0
rect 2628 0 2700 8
rect 2628 8 2700 17
rect 2628 17 2700 26
rect 2628 26 2700 35
rect 2700 -35 2772 -26
rect 2700 -26 2772 -17
rect 2700 -17 2772 -8
rect 2700 -8 2772 0
rect 2700 0 2772 8
rect 2700 8 2772 17
rect 2700 17 2772 26
rect 2700 26 2772 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 2556 316 2628 325
rect 2556 325 2628 334
rect 2556 334 2628 343
rect 2556 343 2628 352
rect 2556 352 2628 360
rect 2556 360 2628 369
rect 2556 369 2628 378
rect 2556 378 2628 387
rect 2628 316 2700 325
rect 2628 325 2700 334
rect 2628 334 2700 343
rect 2628 343 2700 352
rect 2628 352 2700 360
rect 2628 360 2700 369
rect 2628 369 2700 378
rect 2628 378 2700 387
rect 2700 316 2772 325
rect 2700 325 2772 334
rect 2700 334 2772 343
rect 2700 343 2772 352
rect 2700 352 2772 360
rect 2700 360 2772 369
rect 2700 369 2772 378
rect 2700 378 2772 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 2556 668 2628 677
rect 2556 677 2628 686
rect 2556 686 2628 695
rect 2556 695 2628 704
rect 2556 704 2628 712
rect 2556 712 2628 721
rect 2556 721 2628 730
rect 2556 730 2628 739
rect 2628 668 2700 677
rect 2628 677 2700 686
rect 2628 686 2700 695
rect 2628 695 2700 704
rect 2628 704 2700 712
rect 2628 712 2700 721
rect 2628 721 2700 730
rect 2628 730 2700 739
rect 2700 668 2772 677
rect 2700 677 2772 686
rect 2700 686 2772 695
rect 2700 695 2772 704
rect 2700 704 2772 712
rect 2700 712 2772 721
rect 2700 721 2772 730
rect 2700 730 2772 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< v2 >>
rect 2556 -35 2628 -26
rect 2556 -26 2628 -17
rect 2556 -17 2628 -8
rect 2556 -8 2628 0
rect 2556 0 2628 8
rect 2556 8 2628 17
rect 2556 17 2628 26
rect 2556 26 2628 35
rect 2628 -35 2700 -26
rect 2628 -26 2700 -17
rect 2628 -17 2700 -8
rect 2628 -8 2700 0
rect 2628 0 2700 8
rect 2628 8 2700 17
rect 2628 17 2700 26
rect 2628 26 2700 35
rect 2700 -35 2772 -26
rect 2700 -26 2772 -17
rect 2700 -17 2772 -8
rect 2700 -8 2772 0
rect 2700 0 2772 8
rect 2700 8 2772 17
rect 2700 17 2772 26
rect 2700 26 2772 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 2556 316 2628 325
rect 2556 325 2628 334
rect 2556 334 2628 343
rect 2556 343 2628 352
rect 2556 352 2628 360
rect 2556 360 2628 369
rect 2556 369 2628 378
rect 2556 378 2628 387
rect 2628 316 2700 325
rect 2628 325 2700 334
rect 2628 334 2700 343
rect 2628 343 2700 352
rect 2628 352 2700 360
rect 2628 360 2700 369
rect 2628 369 2700 378
rect 2628 378 2700 387
rect 2700 316 2772 325
rect 2700 325 2772 334
rect 2700 334 2772 343
rect 2700 343 2772 352
rect 2700 352 2772 360
rect 2700 360 2772 369
rect 2700 369 2772 378
rect 2700 378 2772 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 2556 668 2628 677
rect 2556 677 2628 686
rect 2556 686 2628 695
rect 2556 695 2628 704
rect 2556 704 2628 712
rect 2556 712 2628 721
rect 2556 721 2628 730
rect 2556 730 2628 739
rect 2628 668 2700 677
rect 2628 677 2700 686
rect 2628 686 2700 695
rect 2628 695 2700 704
rect 2628 704 2700 712
rect 2628 712 2700 721
rect 2628 721 2700 730
rect 2628 730 2700 739
rect 2700 668 2772 677
rect 2700 677 2772 686
rect 2700 686 2772 695
rect 2700 695 2772 704
rect 2700 704 2772 712
rect 2700 712 2772 721
rect 2700 721 2772 730
rect 2700 730 2772 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< viali >>
rect 2556 -35 2628 -26
rect 2556 -26 2628 -17
rect 2556 -17 2628 -8
rect 2556 -8 2628 0
rect 2556 0 2628 8
rect 2556 8 2628 17
rect 2556 17 2628 26
rect 2556 26 2628 35
rect 2628 -35 2700 -26
rect 2628 -26 2700 -17
rect 2628 -17 2700 -8
rect 2628 -8 2700 0
rect 2628 0 2700 8
rect 2628 8 2700 17
rect 2628 17 2700 26
rect 2628 26 2700 35
rect 2700 -35 2772 -26
rect 2700 -26 2772 -17
rect 2700 -17 2772 -8
rect 2700 -8 2772 0
rect 2700 0 2772 8
rect 2700 8 2772 17
rect 2700 17 2772 26
rect 2700 26 2772 35
rect 324 140 396 149
rect 324 149 396 158
rect 324 158 396 167
rect 324 167 396 176
rect 324 176 396 184
rect 324 184 396 193
rect 324 193 396 202
rect 324 202 396 211
rect 396 140 468 149
rect 396 149 468 158
rect 396 158 468 167
rect 396 167 468 176
rect 396 176 468 184
rect 396 184 468 193
rect 396 193 468 202
rect 396 202 468 211
rect 468 140 540 149
rect 468 149 540 158
rect 468 158 540 167
rect 468 167 540 176
rect 468 176 540 184
rect 468 184 540 193
rect 468 193 540 202
rect 468 202 540 211
rect 2556 316 2628 325
rect 2556 325 2628 334
rect 2556 334 2628 343
rect 2556 343 2628 352
rect 2556 352 2628 360
rect 2556 360 2628 369
rect 2556 369 2628 378
rect 2556 378 2628 387
rect 2628 316 2700 325
rect 2628 325 2700 334
rect 2628 334 2700 343
rect 2628 343 2700 352
rect 2628 352 2700 360
rect 2628 360 2700 369
rect 2628 369 2700 378
rect 2628 378 2700 387
rect 2700 316 2772 325
rect 2700 325 2772 334
rect 2700 334 2772 343
rect 2700 343 2772 352
rect 2700 352 2772 360
rect 2700 360 2772 369
rect 2700 369 2772 378
rect 2700 378 2772 387
rect 324 492 396 501
rect 324 501 396 510
rect 324 510 396 519
rect 324 519 396 528
rect 324 528 396 536
rect 324 536 396 545
rect 324 545 396 554
rect 324 554 396 563
rect 396 492 468 501
rect 396 501 468 510
rect 396 510 468 519
rect 396 519 468 528
rect 396 528 468 536
rect 396 536 468 545
rect 396 545 468 554
rect 396 554 468 563
rect 468 492 540 501
rect 468 501 540 510
rect 468 510 540 519
rect 468 519 540 528
rect 468 528 540 536
rect 468 536 540 545
rect 468 545 540 554
rect 468 554 540 563
rect 2556 668 2628 677
rect 2556 677 2628 686
rect 2556 686 2628 695
rect 2556 695 2628 704
rect 2556 704 2628 712
rect 2556 712 2628 721
rect 2556 721 2628 730
rect 2556 730 2628 739
rect 2628 668 2700 677
rect 2628 677 2700 686
rect 2628 686 2700 695
rect 2628 695 2700 704
rect 2628 704 2700 712
rect 2628 712 2700 721
rect 2628 721 2700 730
rect 2628 730 2700 739
rect 2700 668 2772 677
rect 2700 677 2772 686
rect 2700 686 2772 695
rect 2700 695 2772 704
rect 2700 704 2772 712
rect 2700 712 2772 721
rect 2700 721 2772 730
rect 2700 730 2772 739
rect 324 844 396 853
rect 324 853 396 862
rect 324 862 396 871
rect 324 871 396 880
rect 324 880 396 888
rect 324 888 396 897
rect 324 897 396 906
rect 324 906 396 915
rect 396 844 468 853
rect 396 853 468 862
rect 396 862 468 871
rect 396 871 468 880
rect 396 880 468 888
rect 396 888 468 897
rect 396 897 468 906
rect 396 906 468 915
rect 468 844 540 853
rect 468 853 540 862
rect 468 862 540 871
rect 468 871 540 880
rect 468 880 540 888
rect 468 888 540 897
rect 468 897 540 906
rect 468 906 540 915
<< m3 >>
rect 108 -44 2916 44
rect 108 -44 2916 44
rect 2844 44 2916 132
rect 108 132 2556 220
rect 2628 132 2772 220
rect 2844 132 2916 220
rect 108 220 180 308
rect 2844 220 2916 308
rect 108 308 180 396
rect 252 308 324 396
rect 396 308 2916 396
rect 108 396 180 484
rect 2844 396 2916 484
rect 108 484 2772 572
rect 2844 484 2916 572
rect 108 572 180 660
rect 2844 572 2916 660
rect 108 660 180 748
rect 252 660 2916 748
rect 108 748 180 836
rect 108 836 2916 924
rect 108 836 2916 924
<< rm3 >>
rect 2556 132 2628 220
rect 324 308 396 396
<< labels >>
flabel m3 s 108 -44 2916 44 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 108 836 2916 924 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2952 1056
<< end >>
