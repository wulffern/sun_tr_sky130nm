magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 1260 2640
<< locali >>
rect 396 410 564 470
rect 396 1114 564 1174
rect 564 410 624 1174
rect 1152 132 1368 220
rect 288 58 504 118
rect 288 1290 504 1350
rect 720 146 936 206
rect 720 1202 936 1262
rect 288 410 504 470
use SUNTR_PCHDLCM2 M0 
transform 1 0 0 0 1 0
box 0 0 1260 1056
use SUNTR_PCHDLA M1 
transform 1 0 0 0 1 1056
box 0 1056 1260 2640
<< labels >>
flabel locali s 1152 132 1368 220 0 FreeSans 400 0 0 0 B
port 6 nsew signal bidirectional
flabel locali s 288 58 504 118 0 FreeSans 400 0 0 0 S
port 4 nsew signal bidirectional
flabel locali s 288 1290 504 1350 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 720 146 936 206 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 720 1202 936 1262 0 FreeSans 400 0 0 0 CG
port 3 nsew signal bidirectional
flabel locali s 288 410 504 470 0 FreeSans 400 0 0 0 CS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 2640
<< end >>
