magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 2520 1408
<< locali >>
rect 864 234 1032 294
rect 864 938 1032 998
rect 1032 234 1656 294
rect 1032 938 1656 998
rect 1032 234 1092 998
rect 402 146 462 1262
rect 2058 146 2118 1262
rect 834 234 894 470
rect 834 586 894 822
rect 834 938 894 1174
rect 1626 234 1686 470
rect 1626 586 1686 822
rect 1626 938 1686 1174
rect 324 146 540 206
rect 756 234 972 294
<< poly >>
rect 324 158 2196 194
rect 324 510 2196 546
rect 324 862 2196 898
rect 324 1214 2196 1250
<< m2 >>
rect 1656 58 1828 134
rect 1656 586 1828 662
rect 1656 1290 1828 1366
rect 1828 586 2224 662
rect 1828 58 1904 1366
<< m3 >>
rect 2124 586 2324 786
rect 756 0 956 1408
rect 756 0 956 1408
use SUNTR_NCHDL MN0
transform 1 0 0 0 1 0
box 0 0 1260 352
use SUNTR_NCHDL MN1
transform 1 0 0 0 1 352
box 0 352 1260 704
use SUNTR_NCHDL MN2
transform 1 0 0 0 1 704
box 0 704 1260 1056
use SUNTR_NCHDL MN3
transform 1 0 0 0 1 1056
box 0 1056 1260 1408
use SUNTR_PCHDL MP0
transform 1 0 1260 0 1 0
box 1260 0 2520 352
use SUNTR_PCHDL MP1
transform 1 0 1260 0 1 352
box 1260 352 2520 704
use SUNTR_PCHDL MP2
transform 1 0 1260 0 1 704
box 1260 704 2520 1056
use SUNTR_PCHDL MP3
transform 1 0 1260 0 1 1056
box 1260 1056 2520 1408
use SUNTR_cut_M3M4_2x2 xcut0
transform 1 0 2124 0 1 586
box 2124 586 2324 786
use SUNTR_cut_M1M3_2x1 xcut1
transform 1 0 1548 0 1 58
box 1548 58 1748 134
use SUNTR_cut_M1M3_2x1 xcut2
transform 1 0 1548 0 1 586
box 1548 586 1748 662
use SUNTR_cut_M1M3_2x1 xcut3
transform 1 0 1548 0 1 1290
box 1548 1290 1748 1366
use SUNTR_cut_M1M4_2x1 xcut4
transform 1 0 756 0 1 58
box 756 58 956 134
use SUNTR_cut_M1M4_2x1 xcut5
transform 1 0 756 0 1 586
box 756 586 956 662
use SUNTR_cut_M1M4_2x1 xcut6
transform 1 0 756 0 1 762
box 756 762 956 838
use SUNTR_cut_M1M4_2x1 xcut7
transform 1 0 756 0 1 1290
box 756 1290 956 1366
<< labels >>
flabel locali s 324 146 540 206 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 756 234 972 294 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel m3 s 2124 586 2324 786 0 FreeSans 400 0 0 0 VREF
port 3 nsew signal bidirectional
flabel m3 s 756 0 956 1408 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2520 1408
<< end >>
