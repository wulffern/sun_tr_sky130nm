* NGSPICE file created from SUNTR_NCHDL.ext - technology: sky130B

.subckt SUNTR_NCHDL D G S B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=6.156e+11p pd=3.3e+06u as=6.156e+11p ps=3.3e+06u w=1.08e+06u l=180000u
.ends
