magic
tech sky130A
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 2672 4236
<< locali >>
rect 16 16 2656 128
rect 16 16 2656 128
rect 16 16 128 4220
rect 16 4108 2656 4220
rect 2544 16 2656 4220
rect 16 16 2656 128
rect 1480 3438 2056 3658
rect 616 3438 1192 3658
<< ptapc >>
rect 56 32 136 112
rect 136 32 216 112
rect 216 32 296 112
rect 296 32 376 112
rect 376 32 456 112
rect 456 32 536 112
rect 536 32 616 112
rect 616 32 696 112
rect 696 32 776 112
rect 776 32 856 112
rect 856 32 936 112
rect 936 32 1016 112
rect 1016 32 1096 112
rect 1096 32 1176 112
rect 1176 32 1256 112
rect 1256 32 1336 112
rect 1336 32 1416 112
rect 1416 32 1496 112
rect 1496 32 1576 112
rect 1576 32 1656 112
rect 1656 32 1736 112
rect 1736 32 1816 112
rect 1816 32 1896 112
rect 1896 32 1976 112
rect 1976 32 2056 112
rect 2056 32 2136 112
rect 2136 32 2216 112
rect 2216 32 2296 112
rect 2296 32 2376 112
rect 2376 32 2456 112
rect 2456 32 2536 112
rect 2536 32 2616 112
rect 32 38 112 118
rect 32 118 112 198
rect 32 198 112 278
rect 32 278 112 358
rect 32 358 112 438
rect 32 438 112 518
rect 32 518 112 598
rect 32 598 112 678
rect 32 678 112 758
rect 32 758 112 838
rect 32 838 112 918
rect 32 918 112 998
rect 32 998 112 1078
rect 32 1078 112 1158
rect 32 1158 112 1238
rect 32 1238 112 1318
rect 32 1318 112 1398
rect 32 1398 112 1478
rect 32 1478 112 1558
rect 32 1558 112 1638
rect 32 1638 112 1718
rect 32 1718 112 1798
rect 32 1798 112 1878
rect 32 1878 112 1958
rect 32 1958 112 2038
rect 32 2038 112 2118
rect 32 2118 112 2198
rect 32 2198 112 2278
rect 32 2278 112 2358
rect 32 2358 112 2438
rect 32 2438 112 2518
rect 32 2518 112 2598
rect 32 2598 112 2678
rect 32 2678 112 2758
rect 32 2758 112 2838
rect 32 2838 112 2918
rect 32 2918 112 2998
rect 32 2998 112 3078
rect 32 3078 112 3158
rect 32 3158 112 3238
rect 32 3238 112 3318
rect 32 3318 112 3398
rect 32 3398 112 3478
rect 32 3478 112 3558
rect 32 3558 112 3638
rect 32 3638 112 3718
rect 32 3718 112 3798
rect 32 3798 112 3878
rect 32 3878 112 3958
rect 32 3958 112 4038
rect 32 4038 112 4118
rect 32 4118 112 4198
rect 56 4124 136 4204
rect 136 4124 216 4204
rect 216 4124 296 4204
rect 296 4124 376 4204
rect 376 4124 456 4204
rect 456 4124 536 4204
rect 536 4124 616 4204
rect 616 4124 696 4204
rect 696 4124 776 4204
rect 776 4124 856 4204
rect 856 4124 936 4204
rect 936 4124 1016 4204
rect 1016 4124 1096 4204
rect 1096 4124 1176 4204
rect 1176 4124 1256 4204
rect 1256 4124 1336 4204
rect 1336 4124 1416 4204
rect 1416 4124 1496 4204
rect 1496 4124 1576 4204
rect 1576 4124 1656 4204
rect 1656 4124 1736 4204
rect 1736 4124 1816 4204
rect 1816 4124 1896 4204
rect 1896 4124 1976 4204
rect 1976 4124 2056 4204
rect 2056 4124 2136 4204
rect 2136 4124 2216 4204
rect 2216 4124 2296 4204
rect 2296 4124 2376 4204
rect 2376 4124 2456 4204
rect 2456 4124 2536 4204
rect 2536 4124 2616 4204
rect 2560 38 2640 118
rect 2560 118 2640 198
rect 2560 198 2640 278
rect 2560 278 2640 358
rect 2560 358 2640 438
rect 2560 438 2640 518
rect 2560 518 2640 598
rect 2560 598 2640 678
rect 2560 678 2640 758
rect 2560 758 2640 838
rect 2560 838 2640 918
rect 2560 918 2640 998
rect 2560 998 2640 1078
rect 2560 1078 2640 1158
rect 2560 1158 2640 1238
rect 2560 1238 2640 1318
rect 2560 1318 2640 1398
rect 2560 1398 2640 1478
rect 2560 1478 2640 1558
rect 2560 1558 2640 1638
rect 2560 1638 2640 1718
rect 2560 1718 2640 1798
rect 2560 1798 2640 1878
rect 2560 1878 2640 1958
rect 2560 1958 2640 2038
rect 2560 2038 2640 2118
rect 2560 2118 2640 2198
rect 2560 2198 2640 2278
rect 2560 2278 2640 2358
rect 2560 2358 2640 2438
rect 2560 2438 2640 2518
rect 2560 2518 2640 2598
rect 2560 2598 2640 2678
rect 2560 2678 2640 2758
rect 2560 2758 2640 2838
rect 2560 2838 2640 2918
rect 2560 2918 2640 2998
rect 2560 2998 2640 3078
rect 2560 3078 2640 3158
rect 2560 3158 2640 3238
rect 2560 3238 2640 3318
rect 2560 3318 2640 3398
rect 2560 3398 2640 3478
rect 2560 3478 2640 3558
rect 2560 3558 2640 3638
rect 2560 3638 2640 3718
rect 2560 3718 2640 3798
rect 2560 3798 2640 3878
rect 2560 3878 2640 3958
rect 2560 3958 2640 4038
rect 2560 4038 2640 4118
rect 2560 4118 2640 4198
<< ptap >>
rect 0 0 2672 144
rect 0 0 144 4236
rect 0 4092 2672 4236
rect 2528 0 2672 4236
use SUNTR_RES2 XA1
transform 1 0 688 0 1 688
box 688 688 1984 3548
<< labels >>
flabel locali s 16 16 2656 128 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel locali s 1480 3438 2056 3658 0 FreeSans 400 0 0 0 P
port 1 nsew
flabel locali s 616 3438 1192 3658 0 FreeSans 400 0 0 0 N
port 2 nsew
<< end >>
